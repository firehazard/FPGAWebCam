library verilog;
use verilog.vl_types.all;
entity pcpacket_testbench is
end pcpacket_testbench;
