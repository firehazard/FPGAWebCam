library verilog;
use verilog.vl_types.all;
entity edge_detect is
    port(
        clk             : in     vl_logic;
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end edge_detect;
