// Xilinx Verilog netlist produced by netgen application (version G.38)
// Command      : -ofmt verilog -sim temac1.ngd 
// Input file   : temac1.ngd
// Output file  : temac1.v
// Design name  : temac1
// # of Modules : 1
// Xilinx       : C:/Xilinx
// Device       : 2vp20ff896-6

// This verilog netlist is a simulation model and uses simulation 
// primitives which may not represent the true implementation of the 
// device, however the netlist is functionally correct and should not 
// be modified. This file cannot be synthesized and should only be used 
// with supported simulation tools.

`timescale 1 ns/1 ps

module temac1 (
  rxcoreclk, phyemacrxdv, phyemacrxer, emacclienttxretransmit, reset, emacclientrxgoodframe, emacclientrxdvld, emacphytxen, emacphytxer, phyemaccol, 
corehassgmii, clientemacpausereq, phyemaccrs, emacclientrxbadframe, emacclienttxcollision, rxgmiimiiclk, txgmiimiiclk, emacclientrxstatsvld, 
speedis100, emacclienttxstatsvld, speedis10100, clientemactxdvld, txcoreclk, emacclienttxack, clientemactxunderrun, emacclientrxd, 
clientemactxifgdelay, emacclientrxstats, tieemacconfigvec, emacclienttxstats, clientemacpauseval, emacphytxd, clientemactxd, phyemacrxd
);
  input rxcoreclk;
  input phyemacrxdv;
  input phyemacrxer;
  output emacclienttxretransmit;
  input reset;
  output emacclientrxgoodframe;
  output emacclientrxdvld;
  output emacphytxen;
  output emacphytxer;
  input phyemaccol;
  input corehassgmii;
  input clientemacpausereq;
  input phyemaccrs;
  output emacclientrxbadframe;
  output emacclienttxcollision;
  input rxgmiimiiclk;
  input txgmiimiiclk;
  output emacclientrxstatsvld;
  output speedis100;
  output emacclienttxstatsvld;
  output speedis10100;
  input clientemactxdvld;
  input txcoreclk;
  output emacclienttxack;
  input clientemactxunderrun;
  output [7 : 0] emacclientrxd;
  input [7 : 0] clientemactxifgdelay;
  output [26 : 0] emacclientrxstats;
  input [66 : 0] tieemacconfigvec;
  output [31 : 0] emacclienttxstats;
  input [15 : 0] clientemacpauseval;
  output [7 : 0] emacphytxd;
  input [7 : 0] clientemactxd;
  input [7 : 0] phyemacrxd;
  wire N0;
  wire NlwRenamedSig_OI_emacclienttxstatsvld;
  wire NlwRenamedSig_OI_speedis10100;
  wire \NlwRenamedSig_OI_BU2/emacphymclkout ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1/O ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I259/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I272/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I285/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I246/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I233/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I26/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I4/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n004610/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9/O ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1/O ;
  wire \BU2/U0/N66097 ;
  wire \BU2/U0/N66092 ;
  wire \BU2/U0/N66087 ;
  wire \BU2/U0/N66082 ;
  wire \BU2/U0/N66077 ;
  wire \BU2/U0/N66072 ;
  wire \BU2/U0/N66067 ;
  wire \BU2/U0/N66062 ;
  wire \BU2/U0/N66057 ;
  wire \BU2/U0/N66052 ;
  wire \BU2/U0/N66047 ;
  wire \BU2/U0/N66042 ;
  wire \BU2/U0/N66037 ;
  wire \BU2/U0/N66032 ;
  wire \BU2/U0/N66027 ;
  wire \BU2/U0/N65416 ;
  wire \BU2/U0/CHOICE3232 ;
  wire \BU2/U0/N65487 ;
  wire \BU2/U0/N66029 ;
  wire \BU2/U0/CHOICE2804 ;
  wire \BU2/U0/CHOICE3161 ;
  wire \BU2/U0/N61129 ;
  wire \BU2/U0/CHOICE2826 ;
  wire \BU2/U0/CHOICE2844 ;
  wire \BU2/U0/CHOICE2798 ;
  wire \BU2/U0/CHOICE2908 ;
  wire \BU2/U0/CHOICE2633 ;
  wire \BU2/U0/CHOICE2820 ;
  wire \BU2/U0/CHOICE2632 ;
  wire \BU2/U0/CHOICE2981 ;
  wire \BU2/U0/CHOICE3205 ;
  wire \BU2/U0/CHOICE3246 ;
  wire \BU2/U0/CHOICE2793 ;
  wire \BU2/U0/N65464 ;
  wire \BU2/U0/CHOICE3171 ;
  wire \BU2/U0/CHOICE2974 ;
  wire \BU2/U0/CHOICE2929 ;
  wire \BU2/U0/CHOICE3315 ;
  wire \BU2/U0/CHOICE3310 ;
  wire \BU2/U0/N65483 ;
  wire \BU2/U0/CHOICE2815 ;
  wire \BU2/U0/N65440 ;
  wire \BU2/U0/CHOICE2560 ;
  wire \BU2/U0/N66034 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG ;
  wire \BU2/U0/CHOICE2553 ;
  wire \BU2/U0/N66131 ;
  wire \BU2/U0/N66133 ;
  wire \BU2/U0/CHOICE3262 ;
  wire \BU2/U0/CHOICE2846 ;
  wire \BU2/U0/CHOICE2787 ;
  wire \BU2/U0/N65428 ;
  wire \BU2/U0/CHOICE2080 ;
  wire \BU2/U0/N59896 ;
  wire \BU2/U0/CHOICE2079 ;
  wire \BU2/U0/CHOICE2034 ;
  wire \BU2/U0/N65330 ;
  wire \BU2/U0/CHOICE2470 ;
  wire \BU2/U0/CHOICE2031 ;
  wire \BU2/U0/CHOICE2441 ;
  wire \BU2/U0/CHOICE2436 ;
  wire \BU2/U0/CHOICE2027 ;
  wire \BU2/U0/N58329 ;
  wire \BU2/U0/CHOICE2024 ;
  wire \BU2/U0/CHOICE2104 ;
  wire \BU2/U0/CHOICE2020 ;
  wire \BU2/U0/N65448 ;
  wire \BU2/U0/CHOICE2162 ;
  wire \BU2/U0/CHOICE2157 ;
  wire \BU2/U0/CHOICE2277 ;
  wire \BU2/U0/CHOICE2211 ;
  wire \BU2/U0/CHOICE2017 ;
  wire \BU2/U0/N65444 ;
  wire \BU2/U0/N65460 ;
  wire \BU2/U0/N57931 ;
  wire \BU2/U0/CHOICE2013 ;
  wire \BU2/U0/N65456 ;
  wire \BU2/U0/N65764 ;
  wire \BU2/U0/CHOICE2010 ;
  wire \BU2/U0/CHOICE2185 ;
  wire \BU2/U0/CHOICE2152 ;
  wire \BU2/U0/CHOICE2455 ;
  wire \BU2/U0/CHOICE2006 ;
  wire \BU2/U0/CHOICE2126 ;
  wire \BU2/U0/N65412 ;
  wire \BU2/U0/CHOICE2809 ;
  wire \BU2/U0/CHOICE2191 ;
  wire \BU2/U0/N65354 ;
  wire \BU2/U0/CHOICE2516 ;
  wire \BU2/U0/CHOICE2531 ;
  wire \BU2/U0/CHOICE2524 ;
  wire \BU2/U0/CHOICE2003 ;
  wire \BU2/U0/CHOICE2091 ;
  wire \BU2/U0/N65751 ;
  wire \BU2/U0/N50382 ;
  wire \BU2/U0/N50904 ;
  wire \BU2/U0/N66039 ;
  wire \BU2/U0/CHOICE3272 ;
  wire \BU2/U0/N52476 ;
  wire \BU2/U0/CHOICE1677 ;
  wire \BU2/U0/N65792 ;
  wire \BU2/U0/N50348 ;
  wire \BU2/U0/N65808 ;
  wire \BU2/U0/CHOICE1783 ;
  wire \BU2/U0/N66044 ;
  wire \BU2/U0/N65946 ;
  wire \BU2/U0/N50321 ;
  wire \BU2/U0/N51126 ;
  wire \BU2/U0/N52276 ;
  wire \BU2/U0/N65942 ;
  wire \BU2/U0/N51423 ;
  wire \BU2/U0/N65636 ;
  wire \BU2/U0/N65788 ;
  wire \BU2/U0/N50294 ;
  wire \BU2/U0/N50272 ;
  wire \BU2/U0/N65961 ;
  wire \BU2/U0/N65957 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ;
  wire \BU2/U0/N52831 ;
  wire \BU2/U0/N51935 ;
  wire \BU2/U0/N50226 ;
  wire \BU2/U0/N50778 ;
  wire \BU2/U0/N65468 ;
  wire \BU2/U0/CHOICE2849 ;
  wire \BU2/U0/N51052 ;
  wire \BU2/U0/N51594 ;
  wire \BU2/U0/N50196 ;
  wire \BU2/U0/N50568 ;
  wire \BU2/U0/N65648 ;
  wire \BU2/U0/CHOICE2785 ;
  wire \BU2/U0/CHOICE1713 ;
  wire \BU2/U0/N50165 ;
  wire \BU2/U0/N65965 ;
  wire \BU2/U0/N50537 ;
  wire \BU2/U0/N65804 ;
  wire \BU2/U0/N65784 ;
  wire \BU2/U0/CHOICE1874 ;
  wire \BU2/U0/N50134 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0007 ;
  wire \BU2/U0/CHOICE2771 ;
  wire \BU2/U0/CHOICE2768 ;
  wire \BU2/U0/CHOICE1863 ;
  wire \BU2/U0/CHOICE1845 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4366 ;
  wire \BU2/U0/CHOICE2403 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TC_ASSIGN_I0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_C1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4362 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0005 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0007 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0009 ;
  wire \BU2/U0/CHOICE2409 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ;
  wire \BU2/U0/CHOICE2404 ;
  wire \BU2/U0/CHOICE2394 ;
  wire \BU2/U0/N65902 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0011 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0013 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16530 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0008 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0018 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0019 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16535 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0012 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4296 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4290 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo1 ;
  wire \BU2/U0/CHOICE1866 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4299 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4281 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4302 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_N4870 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4284 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_nor_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4287 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0023 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4305 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_37 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_33 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_36 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_32 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_35 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_31 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_34 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_33 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_29 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_32 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt ;
  wire \BU2/U0/N66049 ;
  wire \BU2/U0/CHOICE2628 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4255 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4249 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo21 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4246 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo20 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4243 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo19 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4240 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo18 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4237 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4231 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo16 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4228 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo15 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4225 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4219 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo13 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4216 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo12 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4213 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4207 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo10 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4204 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo9 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4201 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4195 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4192 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4189 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4183 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4180 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4177 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4169 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4166 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4163 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0104 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4234 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo17 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4222 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo14 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0054 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0020 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0023 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0024 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0026 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0027 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0028 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0029 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0030 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0042 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0032 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0033 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0034 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0035 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0036 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0037 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0038 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0039 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0040 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0041 ;
  wire \BU2/U0/CHOICE3132 ;
  wire \BU2/U0/CHOICE3126 ;
  wire \BU2/U0/CHOICE2881 ;
  wire \BU2/U0/CHOICE2870 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0050 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0055 ;
  wire \BU2/U0/N65388 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0062 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0063 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0064 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0096 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0065 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0095 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0066 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0067 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL ;
  wire \BU2/U0/N66187 ;
  wire \BU2/U0/N66054 ;
  wire \BU2/U0/N66195 ;
  wire \BU2/U0/N50513 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_42 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_40 ;
  wire \BU2/U0/N57873 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0110 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_39 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_43 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_46 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_29 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_30 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_37 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_40 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_41 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_42 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_31 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_38 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_41 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_32 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_33 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_34 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_35 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_43 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_36 ;
  wire \BU2/U0/N65780 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0161 ;
  wire \BU2/U0/CHOICE1878 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0175 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0075 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0181 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_36 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0052 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16087 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<9>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<10>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0093 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4210 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo11 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0097 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4198 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo8 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0094 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4186 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0098 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4172 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0103 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4252 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo22 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_45 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_44 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_39 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_35 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_38 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0029 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0030 ;
  wire \BU2/U0/CHOICE1738 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0027 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0044 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0015 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0018 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0021 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0022 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0023 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0024 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0062 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0061 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0060 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0058 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0064 ;
  wire \BU2/U0/CHOICE1831 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0055 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0046 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0059 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0045 ;
  wire \BU2/U0/N66059 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0057 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0056 ;
  wire \BU2/U0/N66064 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0042 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0041 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0040 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0035 ;
  wire \BU2/U0/N65628 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0034 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0043 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0054 ;
  wire \BU2/U0/N65938 ;
  wire \BU2/U0/N54124 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0051 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0050 ;
  wire \BU2/U0/N65934 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0049 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0048 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0047 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0039 ;
  wire \BU2/U0/N65930 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0038 ;
  wire \BU2/U0/N65926 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0037 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0036 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0044 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0053 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0065 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0052 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ;
  wire \BU2/U0/N65776 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_26 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_25 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_24 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI ;
  wire \BU2/U0/N65358 ;
  wire \BU2/U0/CHOICE2486 ;
  wire \BU2/U0/CHOICE2494 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_25 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_23 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_22 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_26 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_30 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_28 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_28 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_24 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_27 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_29 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22745 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV100_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV10_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0063 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_34 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_28 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_27 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0034 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0001 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0000 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CRC1000_EN ;
  wire \BU2/U0/TRIMAC_INST_INT_GMII_RX_DV ;
  wire \BU2/U0/TRIMAC_INST_INT_GMII_RX_ER ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0016 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0017 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0019 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0022 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0023 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0025 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT ;
  wire \BU2/U0/CHOICE2928 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0028 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0029 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0030 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6q ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG5 ;
  wire \BU2/U0/CHOICE2122 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0018 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0024 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT ;
  wire \BU2/U0/CHOICE1868 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WR_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WR_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG5 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0049 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n0006 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG ;
  wire \BU2/U0/CHOICE1120 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_INT_RX_ERR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21520 ;
  wire \BU2/U0/N66216 ;
  wire \BU2/U0/CHOICE3193 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22745 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WR_REG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WR_REG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4378 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0001 ;
  wire \BU2/U0/N66069 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0014 ;
  wire \BU2/U0/N66129 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0044 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4370 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_22 ;
  wire \BU2/U0/N66102 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_INT_RX_DV ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4354 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0000 ;
  wire \BU2/U0/CHOICE1757 ;
  wire \BU2/U0/CHOICE1739 ;
  wire \BU2/U0/CHOICE1725 ;
  wire \BU2/U0/CHOICE1714 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4366 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0016 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4358 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4362 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ;
  wire \BU2/U0/CHOICE3250 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt ;
  wire \BU2/U0/N50978 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5-In ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4354 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_N21825 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0064 ;
  wire \BU2/U0/N66074 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0055 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0046 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0045 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_30 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0057 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0056 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036 ;
  wire \BU2/U0/CHOICE2587 ;
  wire \BU2/U0/N65432 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0042 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0041 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0040 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0035 ;
  wire \BU2/U0/N65906 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0034 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0043 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0054 ;
  wire \BU2/U0/N65922 ;
  wire \BU2/U0/N66079 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0051 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0050 ;
  wire \BU2/U0/N65918 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0049 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0048 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0047 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0039 ;
  wire \BU2/U0/N65914 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0038 ;
  wire \BU2/U0/N65910 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0037 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0036 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0044 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0053 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0065 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0052 ;
  wire \BU2/U0/N65772 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4335 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4331 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4327 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4323 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4319 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4315 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>_cyo ;
  wire \BU2/U0/N52548 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3 ;
  wire \BU2/U0/CHOICE2595 ;
  wire \BU2/U0/CHOICE2590 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4339 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4343 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026 ;
  wire \BU2/U0/N50462 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22904 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG ;
  wire \BU2/U0/N66231 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0058 ;
  wire \BU2/U0/N53888 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010 ;
  wire \BU2/U0/CHOICE3208 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21559 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n0000 ;
  wire \BU2/U0/N65436 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ;
  wire \BU2/U0/CHOICE2701 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4622 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4619 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4616 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4613 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4610 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4607 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4604 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4596 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4592 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4588 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[15] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[14] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4566 ;
  wire \BU2/U0/CHOICE3153 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4562 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[6] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[5] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4548 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt ;
  wire \BU2/U0/CHOICE2918 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4542 ;
  wire \BU2/U0/CHOICE3115 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4534 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4530 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4526 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4522 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4518 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_27 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4514 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4510 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_23 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[5] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4506 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_25 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[3] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4502 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4498 ;
  wire \BU2/U0/N65392 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[4] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[13] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4494 ;
  wire \BU2/U0/CHOICE1830 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4490 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4486 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4482 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4478 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4474 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4470 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0084 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH ;
  wire \BU2/U0/N66255 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4446 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4438 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4434 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4430 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4426 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4422 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4418 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4414 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4410 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4406 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4402 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4398 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4394 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4390 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0144 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0132 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0131 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0130 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0129 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0128 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0512 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0511 ;
  wire \BU2/U0/N66193 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0475 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0179 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0463 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0462 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0461 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0460 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0459 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0350 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458 ;
  wire \BU2/U0/N66185 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0171 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD ;
  wire \BU2/U0/N66126 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0447 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0446 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0291 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0445 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0287 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0038 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[9] ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0082 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0104 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0081 ;
  wire \BU2/U0/CHOICE3268 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0060 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0111 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[18] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0068 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0080 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0123 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt ;
  wire \BU2/U0/CHOICE2087 ;
  wire \BU2/U0/CHOICE2216 ;
  wire \BU2/U0/CHOICE2209 ;
  wire \BU2/U0/N65984 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0076 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_CONTROL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0074 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0191 ;
  wire \BU2/U0/N53396 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21490 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0146 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0079 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0115 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0078 ;
  wire \BU2/U0/N51861 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0086 ;
  wire \BU2/U0/N66253 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_39 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt ;
  wire \BU2/U0/N52182 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0070 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0102 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[10] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0165 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG ;
  wire \BU2/U0/CHOICE2237 ;
  wire \BU2/U0/CHOICE2230 ;
  wire \BU2/U0/CHOICE2250 ;
  wire \BU2/U0/CHOICE2243 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0061 ;
  wire \BU2/U0/N66250 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0174 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0060 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16128 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0095 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0186 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_43 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0188 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0189 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0063 ;
  wire \BU2/U0/N65592 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0196 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0192 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0058 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_24 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0200 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0202 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0057 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0198 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ;
  wire \BU2/U0/CHOICE2540 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22904 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_65 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_60 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0056 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_62 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_49 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_DONE ;
  wire \BU2/U0/N65420 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012 ;
  wire \BU2/U0/CHOICE2940 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_46 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_50 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0319 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_64 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_47 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_51 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_47 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0047 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0092 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_48 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_52 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_48 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0046 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_53 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_49 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11 ;
  wire \BU2/U0/N65882 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[2] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0449 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_45 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0302 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_56 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[17] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21290 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[16] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_46 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_45 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0045 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_59 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_64 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64 ;
  wire \BU2/U0/CHOICE2048 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_60 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[15] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[13] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_50 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_55 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_50 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[14] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN__n0033 ;
  wire \BU2/U0/N65452 ;
  wire \BU2/U0/CHOICE2117 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[12] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_51 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_51 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_56 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[11] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_52 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_52 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_57 ;
  wire \BU2/U0/CHOICE3145 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ;
  wire \BU2/U0/CHOICE3141 ;
  wire \BU2/U0/CHOICE3136 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_53 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_58 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_53 ;
  wire \BU2/U0/CHOICE3182 ;
  wire \BU2/U0/CHOICE3181 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0077 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_54 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_59 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_54 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_55 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_60 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_55 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0077 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0177 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8 ;
  wire \BU2/U0/N65396 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[3] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[12] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_56 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_61 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_57 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_62 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_57 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1 ;
  wire \BU2/U0/CHOICE2778 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_64 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[5] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_59 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_58 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_63 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_58 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[6] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[7] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_67 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[8] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_62 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_61 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_66 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_61 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0218 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0153 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_63 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_69 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_63 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_68 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_49 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_44 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_48 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_44 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_45 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_46 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0443 ;
  wire \BU2/U0/CHOICE3129 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ;
  wire \BU2/U0/N66084 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0450 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0167 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0451 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0308 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0452 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0313 ;
  wire \BU2/U0/CHOICE2709 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ;
  wire \BU2/U0/N50430 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0456 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0457 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0173 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1 ;
  wire \BU2/U0/CHOICE1790 ;
  wire \BU2/U0/N66089 ;
  wire \BU2/U0/CHOICE3286 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022__n0002 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0464 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DELAYED ;
  wire \BU2/U0/N65254 ;
  wire \BU2/U0/CHOICE3329 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0531 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ;
  wire \BU2/U0/N50821 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ;
  wire \BU2/U0/N51266 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0062 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0471 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0472 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0473 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0273 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0474 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ;
  wire \BU2/U0/N65408 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0510 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[1] ;
  wire \BU2/U0/N65400 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[2] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[11] ;
  wire \BU2/U0/N66094 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0514 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0513 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0523 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0524 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0525 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4600 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0527 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0528 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4538 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0530 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0226 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4625 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0061 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4442 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0022 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ;
  wire \BU2/U0/N51500 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197 ;
  wire \BU2/U0/N66288 ;
  wire \BU2/U0/N53310 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ;
  wire \BU2/U0/N52675 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<8>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<9>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ;
  wire \BU2/U0/N66290 ;
  wire \BU2/U0/N53474 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1__n0000 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_N17122 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>__net3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[0] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TC ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TC ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TC ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TC ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TC_ASSIGN_I0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ0 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_C1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_24 ;
  wire \BU2/U0/N52594 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_26 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_23 ;
  wire \BU2/U0/CHOICE1820 ;
  wire \BU2/U0/CHOICE1819 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_25 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_22 ;
  wire \BU2/U0/N66295 ;
  wire \BU2/U0/N53520 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_24 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0068 ;
  wire \BU2/U0/N53563 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[5] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_25 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_23 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_22 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[3] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_26 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_26 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_30 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_28 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_28 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_24 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_27 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_29 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_27 ;
  wire \BU2/U0/CHOICE2389 ;
  wire \BU2/U0/N65472 ;
  wire \BU2/U0/CHOICE2384 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[8] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[17] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4152 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4148 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4144 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4140 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4136 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4132 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4128 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4124 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4120 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4116 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4112 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ;
  wire \BU2/U0/N65404 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[1] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[10] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1 ;
  wire \BU2/U0/N51803 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16092 ;
  wire \BU2/U0/N65280 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[7] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[16] ;
  wire \BU2/U0/CHOICE1809 ;
  wire \BU2/U0/CHOICE1804 ;
  wire \BU2/U0/CHOICE1791 ;
  wire \BU2/U0/CHOICE1844 ;
  wire \BU2/U0/N56896 ;
  wire \BU2/U0/CHOICE1703 ;
  wire \BU2/U0/CHOICE1698 ;
  wire \BU2/U0/CHOICE1685 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In ;
  wire \BU2/U0/CHOICE1684 ;
  wire \BU2/U0/N65284 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ;
  wire \BU2/U0/N66312 ;
  wire \BU2/U0/N65067 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4156 ;
  wire \BU2/U0/CHOICE3085 ;
  wire \BU2/U0/CHOICE3082 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0001 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_28 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_25 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_27 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[14] ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0060 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TC ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4q ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ;
  wire \BU2/U0/CHOICE2726 ;
  wire \BU2/U0/CHOICE2752 ;
  wire \BU2/U0/CHOICE2720 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_TX_EN_DELAY ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0011 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0012 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0014 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0016 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0017 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0018 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0020 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_CRS ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0022 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0013 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES_PRE_REG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0019 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ;
  wire \BU2/U0/TRIMAC_INST_TXGEN__n0034 ;
  wire \BU2/U0/CHOICE1945 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In ;
  wire \BU2/U0/CHOICE2177 ;
  wire \BU2/U0/CHOICE2173 ;
  wire \BU2/U0/CHOICE2833 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0012 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0066 ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_ACK_EARLY_IN ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_ACK_IN ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19418 ;
  wire \BU2/U0/N66190 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ;
  wire \BU2/U0/CHOICE3332 ;
  wire \BU2/U0/N65986 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ;
  wire \BU2/U0/N61770 ;
  wire \BU2/U0/CHOICE2706 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ;
  wire \BU2/U0/CHOICE2693 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ;
  wire \BU2/U0/CHOICE2702 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ;
  wire \BU2/U0/N66135 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ;
  wire \BU2/U0/N66317 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ;
  wire \BU2/U0/CHOICE2085 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD ;
  wire \BU2/U0/N65368 ;
  wire \BU2/U0/CHOICE3073 ;
  wire \BU2/U0/CHOICE3067 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ;
  wire \BU2/U0/CHOICE1339 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354 ;
  wire \BU2/U0/N62536 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0022 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0454 ;
  wire \BU2/U0/CHOICE2651 ;
  wire \BU2/U0/N66248 ;
  wire \BU2/U0/CHOICE3109 ;
  wire \BU2/U0/CHOICE3106 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0011 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_COMB ;
  wire \BU2/U0/CHOICE2949 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ;
  wire \BU2/U0/N66297 ;
  wire \BU2/U0/N66180 ;
  wire \BU2/U0/N65372 ;
  wire \BU2/U0/CHOICE3097 ;
  wire \BU2/U0/CHOICE3091 ;
  wire \BU2/U0/CHOICE3061 ;
  wire \BU2/U0/CHOICE3058 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0015 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0069 ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_UNDERRUN_OUT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0004 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0007 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0008 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0009 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0010 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0011 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT ;
  wire \BU2/U0/CHOICE2463 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ;
  wire \BU2/U0/N59033 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0012 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0013 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0014 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0038 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0039 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0021 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_N18510 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0051 ;
  wire \BU2/U0/CHOICE2201 ;
  wire \BU2/U0/CHOICE2197 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_21 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_22 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_20 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_21 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_19 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_20 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_18 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_17 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_19 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_17 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_18 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_16 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_17 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_15 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_16 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_14 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_15 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_13 ;
  wire \BU2/U0/CHOICE3259 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_14 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_12 ;
  wire \BU2/U0/N65350 ;
  wire \BU2/U0/CHOICE2716 ;
  wire \BU2/U0/CHOICE2730 ;
  wire \BU2/U0/CHOICE2735 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_13 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_11 ;
  wire \BU2/U0/N65376 ;
  wire \BU2/U0/CHOICE3050 ;
  wire \BU2/U0/CHOICE3044 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_12 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_10 ;
  wire \BU2/U0/CHOICE2839 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_11 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_9 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_10 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_8 ;
  wire \BU2/U0/N65743 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_9 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_7 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 ;
  wire \BU2/U0/N66330 ;
  wire \BU2/U0/CHOICE2680 ;
  wire \BU2/U0/CHOICE2673 ;
  wire \BU2/U0/N65878 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_6 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_8 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_6 ;
  wire \BU2/U0/N65747 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_7 ;
  wire \BU2/U0/N66116 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_21 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_20 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_5 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_18 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_42 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_5 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_4 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_41 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_3 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_4 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_40 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_2 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_3 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_2 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_2 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_38 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_0 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_0 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_37 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_0 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_5 ;
  wire \BU2/U0/CHOICE2600 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0008 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_13 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_12 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG ;
  wire \BU2/U0/CHOICE2501 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_9 ;
  wire \BU2/U0/CHOICE2049 ;
  wire \BU2/U0/CHOICE2041 ;
  wire \BU2/U0/CHOICE2038 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_10 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_14 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_15 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_11 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_16 ;
  wire \BU2/U0/N60912 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0011 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_19 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0021 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0014 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_END_OF_TX ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_8 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0022 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0007 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_4 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX ;
  wire \BU2/U0/TRIMAC_INST_FLOW_PAUSE_REQ_LOCAL ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE__n0000 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_COMB ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_COMB ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_7 ;
  wire \BU2/U0/N52009 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4358 ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_VLAN_ENABLE_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0059 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL ;
  wire \BU2/U0/TRIMAC_INST_FLOW__n0007 ;
  wire \BU2/U0/TRIMAC_INST_FLOW__n0001 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ;
  wire \BU2/U0/TRIMAC_INST_FLOW__n0002 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ;
  wire \BU2/U0/TRIMAC_INST_FLOW__n0003 ;
  wire \BU2/U0/CHOICE2900 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ;
  wire \BU2/U0/CHOICE2899 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014 ;
  wire \BU2/U0/TRIMAC_INST_INT_EXTENSION ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1 ;
  wire \BU2/U0/N53281 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ;
  wire \BU2/U0/N65588 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0059 ;
  wire \BU2/U0/N65768 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In ;
  wire \BU2/U0/CHOICE2994 ;
  wire \BU2/U0/N65873 ;
  wire \BU2/U0/CHOICE2857 ;
  wire \BU2/U0/CHOICE2867 ;
  wire \BU2/U0/CHOICE2863 ;
  wire \BU2/U0/CHOICE3015 ;
  wire \BU2/U0/CHOICE3012 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In ;
  wire \BU2/U0/CHOICE2688 ;
  wire \BU2/U0/N65424 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0046 ;
  wire \BU2/U0/N65527 ;
  wire \BU2/U0/CHOICE3237 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022__n0002 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ;
  wire \BU2/U0/CHOICE3038 ;
  wire \BU2/U0/CHOICE3035 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0016 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ;
  wire \BU2/U0/N66138 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD ;
  wire \BU2/U0/N65380 ;
  wire \BU2/U0/CHOICE3004 ;
  wire \BU2/U0/CHOICE2998 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_26 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC ;
  wire \BU2/U0/N65384 ;
  wire \BU2/U0/CHOICE3027 ;
  wire \BU2/U0/CHOICE3021 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4293 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ;
  wire \BU2/U0/CHOICE2987 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_CONTROL_COMPLETE ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ;
  wire \BU2/U0/N65476 ;
  wire \BU2/U0/N65478 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_N17850 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ;
  wire \BU2/U0/N66099 ;
  wire \BU2/U0/CHOICE2875 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 ;
  wire \BU2/U0/CHOICE2262 ;
  wire \BU2/U0/CHOICE2257 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0011 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0012 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0054 ;
  wire \BU2/U0/CHOICE3280 ;
  wire \BU2/U0/CHOICE2045 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt ;
  wire \BU2/U0/N65759 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_WR_EN ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0453 ;
  wire \BU2/U0/CHOICE2430 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0315 ;
  wire \BU2/U0/CHOICE2424 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0020 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ;
  wire \BU2/U0/CHOICE2655 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0014 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_N4073 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0526 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0016 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4378 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4370 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ;
  wire \BU2/U0/N65520 ;
  wire \BU2/U0/CHOICE2373 ;
  wire \BU2/U0/N65516 ;
  wire \BU2/U0/CHOICE2349 ;
  wire \BU2/U0/N65512 ;
  wire \BU2/U0/CHOICE2361 ;
  wire \BU2/U0/N65508 ;
  wire \BU2/U0/CHOICE2337 ;
  wire \BU2/U0/N65504 ;
  wire \BU2/U0/CHOICE2313 ;
  wire \BU2/U0/N65500 ;
  wire \BU2/U0/CHOICE2325 ;
  wire \BU2/U0/N65496 ;
  wire \BU2/U0/CHOICE2301 ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_INT_ALIGNMENT_ERR_PULSE ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2 ;
  wire \BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2 ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4374 ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4374 ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_N18517 ;
  wire \BU2/U0/N65492 ;
  wire \BU2/U0/CHOICE2289 ;
  wire \BU2/U0/CHOICE1724 ;
  wire \BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ;
  wire \BU2/U0/N66008 ;
  wire \BU2/U0/CHOICE1379 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX__n0067 ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ;
  wire \BU2/U0/address_valid_early ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/CE ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/CE ;
  wire GSR = glbl.GSR;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_CRS.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1.GSR.OR ;
  wire \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2.GSR.OR ;
  wire NLW_VCC_O_UNCONNECTED;
  wire GND;
  wire VCC;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[4]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[5]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[6]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[7]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[8]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[9]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[10]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[11]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[12]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[13]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[14]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[15]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[16]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[17]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[18]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[19]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[20]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[21]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[22]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[23]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[24]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[25]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[26]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[27]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[28]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[29]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[30]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[31]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[11]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[12]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[13]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[14]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[15]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[16]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[17]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[18]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[19]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[20]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[21]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[22]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[23]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[24]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[25]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[26]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[27]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[28]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[29]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[30]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[31]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[4]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[5]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[6]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[7]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[8]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[9]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[10]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[11]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[12]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[13]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[14]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[15]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[16]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[17]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[18]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[19]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[20]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[21]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[22]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[23]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[24]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[25]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[26]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[27]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[28]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[29]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[30]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[31]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[11]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[12]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[13]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[14]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[15]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[16]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[17]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[18]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[19]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[20]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[21]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[22]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[23]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[24]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[25]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[26]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[27]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[28]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[29]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[30]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[31]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[0]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[1]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[2]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[3]_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REGPREDELGEN_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_srl_0_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_TXGEN_BYTECNTSRL_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_FLOW_TX_MUX_ACK_OUT2_O_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/SRL16E_Q15_UNCONNECTED ;
  wire \NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/SRL16E_Q15_UNCONNECTED ;
  wire [7 : 0] emacphytxd_0;
  wire [7 : 0] phyemacrxd_1;
  wire [7 : 0] clientemactxd_2;
  wire [7 : 0] clientemactxifgdelay_3;
  wire [15 : 0] clientemacpauseval_4;
  wire [7 : 0] emacclientrxd_5;
  wire [26 : 2] emacclientrxstats_6;
  wire [1 : 0] NlwRenamedSig_OI_emacclientrxstats;
  wire [66 : 0] tieemacconfigvec_7;
  wire [2 : 1] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q ;
  wire [10 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER ;
  wire [10 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE ;
  wire [5 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE ;
  wire [10 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 ;
  wire [5 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH ;
  wire [5 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH ;
  wire [5 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0296 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0299 ;
  wire [31 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0297 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0116_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0114_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0113_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0112_Xo ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0317 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0101_Xo ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 ;
  wire [3 : 3] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0118_Xo ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0318 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo ;
  wire [47 : 0] \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 ;
  wire [13 : 0] \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_INT_RXD ;
  wire [15 : 8] \BU2/U0/TRIMAC_INST_RXGEN__n0109 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RXD_ALIGNMENT_ERR_RD ;
  wire [8 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR ;
  wire [8 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0297 ;
  wire [31 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo ;
  wire [9 : 1] \BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0116_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0114_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0113_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0112_Xo ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0277 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0277 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0101_Xo ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0294 ;
  wire [3 : 3] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0118_Xo ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0318 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0317 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo ;
  wire [8 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 ;
  wire [8 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 ;
  wire [18 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 ;
  wire [18 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT ;
  wire [15 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN ;
  wire [8 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC ;
  wire [2 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY ;
  wire [9 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT ;
  wire [14 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC ;
  wire [18 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 ;
  wire [9 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 ;
  wire [14 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 ;
  wire [13 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE ;
  wire [7 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED ;
  wire [7 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0299 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 ;
  wire [7 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS ;
  wire [3 : 3] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0100 ;
  wire [9 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN__n0106 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN__n0108 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST ;
  wire [13 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY ;
  wire [9 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 ;
  wire [2 : 2] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0296 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE ;
  wire [6 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT ;
  wire [12 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 ;
  wire [12 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 ;
  wire [12 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR ;
  wire [15 : 0] \BU2/U0/TRIMAC_INST_TXGEN__n0035 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN__n0037 ;
  wire [1 : 0] \BU2/U0/TRIMAC_INST_TXGEN__n0038 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_TXGEN__n0039 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX__n0014 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL ;
  wire [15 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD ;
  wire [4 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 ;
  wire [47 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n0007 ;
  wire [4 : 0] \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY ;
  wire [4 : 0] \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT ;
  wire [15 : 6] \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT ;
  wire [5 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA ;
  wire [4 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT ;
  wire [15 : 0] \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX ;
  wire [15 : 0] \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_RXGEN_DATA ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST__n0009 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 ;
  wire [11 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST__n0012 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST__n0011 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 ;
  wire [3 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002 ;
  wire [0 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY ;
  wire [2 : 0] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY ;
  wire [1 : 1] \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002 ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY ;
  wire [7 : 0] \BU2/U0/TRIMAC_INST_INT_GMII_RXD ;
  assign
    emacclientrxd[7] = emacclientrxd_5[7],
    emacclientrxd[6] = emacclientrxd_5[6],
    emacclientrxd[5] = emacclientrxd_5[5],
    emacclientrxd[4] = emacclientrxd_5[4],
    emacclientrxd[3] = emacclientrxd_5[3],
    emacclientrxd[2] = emacclientrxd_5[2],
    emacclientrxd[1] = emacclientrxd_5[1],
    emacclientrxd[0] = emacclientrxd_5[0],
    clientemactxifgdelay_3[7] = clientemactxifgdelay[7],
    clientemactxifgdelay_3[6] = clientemactxifgdelay[6],
    clientemactxifgdelay_3[5] = clientemactxifgdelay[5],
    clientemactxifgdelay_3[4] = clientemactxifgdelay[4],
    clientemactxifgdelay_3[3] = clientemactxifgdelay[3],
    clientemactxifgdelay_3[2] = clientemactxifgdelay[2],
    clientemactxifgdelay_3[1] = clientemactxifgdelay[1],
    clientemactxifgdelay_3[0] = clientemactxifgdelay[0],
    emacclientrxstats[26] = emacclientrxstats_6[26],
    emacclientrxstats[25] = emacclientrxstats_6[25],
    emacclientrxstats[24] = emacclientrxstats_6[24],
    emacclientrxstats[23] = emacclientrxstats_6[23],
    emacclientrxstats[22] = emacclientrxstats_6[22],
    emacclientrxstats[21] = emacclientrxstats_6[21],
    emacclientrxstats[20] = emacclientrxstats_6[20],
    emacclientrxstats[19] = emacclientrxstats_6[19],
    emacclientrxstats[18] = emacclientrxstats_6[18],
    emacclientrxstats[17] = emacclientrxstats_6[17],
    emacclientrxstats[16] = emacclientrxstats_6[16],
    emacclientrxstats[15] = emacclientrxstats_6[15],
    emacclientrxstats[14] = emacclientrxstats_6[14],
    emacclientrxstats[13] = emacclientrxstats_6[13],
    emacclientrxstats[12] = emacclientrxstats_6[12],
    emacclientrxstats[11] = emacclientrxstats_6[11],
    emacclientrxstats[10] = emacclientrxstats_6[10],
    emacclientrxstats[9] = emacclientrxstats_6[9],
    emacclientrxstats[8] = emacclientrxstats_6[8],
    emacclientrxstats[7] = emacclientrxstats_6[7],
    emacclientrxstats[6] = emacclientrxstats_6[6],
    emacclientrxstats[5] = emacclientrxstats_6[5],
    emacclientrxstats[4] = emacclientrxstats_6[4],
    emacclientrxstats[3] = emacclientrxstats_6[3],
    emacclientrxstats[2] = emacclientrxstats_6[2],
    emacclientrxstats[1] = NlwRenamedSig_OI_emacclientrxstats[1],
    emacclientrxstats[0] = NlwRenamedSig_OI_emacclientrxstats[0],
    tieemacconfigvec_7[66] = tieemacconfigvec[66],
    tieemacconfigvec_7[65] = tieemacconfigvec[65],
    tieemacconfigvec_7[64] = tieemacconfigvec[64],
    tieemacconfigvec_7[63] = tieemacconfigvec[63],
    tieemacconfigvec_7[62] = tieemacconfigvec[62],
    tieemacconfigvec_7[61] = tieemacconfigvec[61],
    tieemacconfigvec_7[60] = tieemacconfigvec[60],
    tieemacconfigvec_7[59] = tieemacconfigvec[59],
    tieemacconfigvec_7[58] = tieemacconfigvec[58],
    tieemacconfigvec_7[57] = tieemacconfigvec[57],
    tieemacconfigvec_7[56] = tieemacconfigvec[56],
    tieemacconfigvec_7[55] = tieemacconfigvec[55],
    tieemacconfigvec_7[54] = tieemacconfigvec[54],
    tieemacconfigvec_7[53] = tieemacconfigvec[53],
    tieemacconfigvec_7[52] = tieemacconfigvec[52],
    tieemacconfigvec_7[51] = tieemacconfigvec[51],
    tieemacconfigvec_7[50] = tieemacconfigvec[50],
    tieemacconfigvec_7[49] = tieemacconfigvec[49],
    tieemacconfigvec_7[48] = tieemacconfigvec[48],
    tieemacconfigvec_7[47] = tieemacconfigvec[47],
    tieemacconfigvec_7[46] = tieemacconfigvec[46],
    tieemacconfigvec_7[45] = tieemacconfigvec[45],
    tieemacconfigvec_7[44] = tieemacconfigvec[44],
    tieemacconfigvec_7[43] = tieemacconfigvec[43],
    tieemacconfigvec_7[42] = tieemacconfigvec[42],
    tieemacconfigvec_7[41] = tieemacconfigvec[41],
    tieemacconfigvec_7[40] = tieemacconfigvec[40],
    tieemacconfigvec_7[39] = tieemacconfigvec[39],
    tieemacconfigvec_7[38] = tieemacconfigvec[38],
    tieemacconfigvec_7[37] = tieemacconfigvec[37],
    tieemacconfigvec_7[36] = tieemacconfigvec[36],
    tieemacconfigvec_7[35] = tieemacconfigvec[35],
    tieemacconfigvec_7[34] = tieemacconfigvec[34],
    tieemacconfigvec_7[33] = tieemacconfigvec[33],
    tieemacconfigvec_7[32] = tieemacconfigvec[32],
    tieemacconfigvec_7[31] = tieemacconfigvec[31],
    tieemacconfigvec_7[30] = tieemacconfigvec[30],
    tieemacconfigvec_7[29] = tieemacconfigvec[29],
    tieemacconfigvec_7[28] = tieemacconfigvec[28],
    tieemacconfigvec_7[27] = tieemacconfigvec[27],
    tieemacconfigvec_7[26] = tieemacconfigvec[26],
    tieemacconfigvec_7[25] = tieemacconfigvec[25],
    tieemacconfigvec_7[24] = tieemacconfigvec[24],
    tieemacconfigvec_7[23] = tieemacconfigvec[23],
    tieemacconfigvec_7[22] = tieemacconfigvec[22],
    tieemacconfigvec_7[21] = tieemacconfigvec[21],
    tieemacconfigvec_7[20] = tieemacconfigvec[20],
    tieemacconfigvec_7[19] = tieemacconfigvec[19],
    tieemacconfigvec_7[18] = tieemacconfigvec[18],
    tieemacconfigvec_7[17] = tieemacconfigvec[17],
    tieemacconfigvec_7[16] = tieemacconfigvec[16],
    tieemacconfigvec_7[15] = tieemacconfigvec[15],
    tieemacconfigvec_7[14] = tieemacconfigvec[14],
    tieemacconfigvec_7[13] = tieemacconfigvec[13],
    tieemacconfigvec_7[12] = tieemacconfigvec[12],
    tieemacconfigvec_7[11] = tieemacconfigvec[11],
    tieemacconfigvec_7[10] = tieemacconfigvec[10],
    tieemacconfigvec_7[9] = tieemacconfigvec[9],
    tieemacconfigvec_7[8] = tieemacconfigvec[8],
    tieemacconfigvec_7[7] = tieemacconfigvec[7],
    tieemacconfigvec_7[6] = tieemacconfigvec[6],
    tieemacconfigvec_7[5] = tieemacconfigvec[5],
    tieemacconfigvec_7[4] = tieemacconfigvec[4],
    tieemacconfigvec_7[3] = tieemacconfigvec[3],
    tieemacconfigvec_7[2] = tieemacconfigvec[2],
    tieemacconfigvec_7[1] = tieemacconfigvec[1],
    tieemacconfigvec_7[0] = tieemacconfigvec[0],
    emacclienttxstats[29] = \NlwRenamedSig_OI_BU2/emacphymclkout ,
    emacclienttxstats[24] = \NlwRenamedSig_OI_BU2/emacphymclkout ,
    clientemacpauseval_4[15] = clientemacpauseval[15],
    clientemacpauseval_4[14] = clientemacpauseval[14],
    clientemacpauseval_4[13] = clientemacpauseval[13],
    clientemacpauseval_4[12] = clientemacpauseval[12],
    clientemacpauseval_4[11] = clientemacpauseval[11],
    clientemacpauseval_4[10] = clientemacpauseval[10],
    clientemacpauseval_4[9] = clientemacpauseval[9],
    clientemacpauseval_4[8] = clientemacpauseval[8],
    clientemacpauseval_4[7] = clientemacpauseval[7],
    clientemacpauseval_4[6] = clientemacpauseval[6],
    clientemacpauseval_4[5] = clientemacpauseval[5],
    clientemacpauseval_4[4] = clientemacpauseval[4],
    clientemacpauseval_4[3] = clientemacpauseval[3],
    clientemacpauseval_4[2] = clientemacpauseval[2],
    clientemacpauseval_4[1] = clientemacpauseval[1],
    clientemacpauseval_4[0] = clientemacpauseval[0],
    emacphytxd[7] = emacphytxd_0[7],
    emacphytxd[6] = emacphytxd_0[6],
    emacphytxd[5] = emacphytxd_0[5],
    emacphytxd[4] = emacphytxd_0[4],
    emacphytxd[3] = emacphytxd_0[3],
    emacphytxd[2] = emacphytxd_0[2],
    emacphytxd[1] = emacphytxd_0[1],
    emacphytxd[0] = emacphytxd_0[0],
    clientemactxd_2[7] = clientemactxd[7],
    clientemactxd_2[6] = clientemactxd[6],
    clientemactxd_2[5] = clientemactxd[5],
    clientemactxd_2[4] = clientemactxd[4],
    clientemactxd_2[3] = clientemactxd[3],
    clientemactxd_2[2] = clientemactxd[2],
    clientemactxd_2[1] = clientemactxd[1],
    clientemactxd_2[0] = clientemactxd[0],
    phyemacrxd_1[7] = phyemacrxd[7],
    phyemacrxd_1[6] = phyemacrxd[6],
    phyemacrxd_1[5] = phyemacrxd[5],
    phyemacrxd_1[4] = phyemacrxd[4],
    phyemacrxd_1[3] = phyemacrxd[3],
    phyemacrxd_1[2] = phyemacrxd[2],
    phyemacrxd_1[1] = phyemacrxd[1],
    phyemacrxd_1[0] = phyemacrxd[0],
    emacclienttxstatsvld = NlwRenamedSig_OI_emacclienttxstatsvld,
    speedis10100 = NlwRenamedSig_OI_speedis10100;
  X_ONE VCC_8 (
    .O(NLW_VCC_O_UNCONNECTED)
  );
  X_ZERO GND_9 (
    .O(N0)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n000515 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n000515  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC ),
    .ADR1(\BU2/U0/CHOICE3329 ),
    .ADR2(\BU2/U0/CHOICE3332 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n000515/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .O(\BU2/U0/N66102 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<7>1/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/CHOICE2787 ),
    .ADR2(\BU2/U0/CHOICE2793 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>38/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/CHOICE2798 ),
    .ADR2(\BU2/U0/CHOICE2804 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>38/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117 .INIT = 16'hF200;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_EXTENSION ),
    .ADR2(\BU2/U0/CHOICE1868 ),
    .ADR3(\BU2/U0/CHOICE1866 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW117/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117 .INIT = 16'hFF8A;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117  (
    .ADR0(\BU2/U0/CHOICE1878 ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_EXTENSION ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .ADR3(\BU2/U0/CHOICE1874 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW117/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/CHOICE2820 ),
    .ADR2(\BU2/U0/CHOICE2826 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>38/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/CHOICE2809 ),
    .ADR2(\BU2/U0/CHOICE2815 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>38/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<4>1/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<5>1/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<6>1/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM1/O ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[15] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[6] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16_SW0/O ),
    .O(\BU2/U0/N65284 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00021 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00021  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00021/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .O(\BU2/U0/N66116 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61  (
    .ADR0(\BU2/U0/N66116 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_61/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_6 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [7]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_71/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_7 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [8]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_81/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_8 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [9]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_91/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_9 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [10]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_101/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_10 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [11]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_111/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_11 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [12]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_121/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_12 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [13]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_131/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_13 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_AVAIL_OUT_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_AVAIL_OUT_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_AVAIL_OUT_Result1/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .O(\BU2/U0/N66126 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424_10 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424_10  (
    .ADR0(\BU2/U0/N53281 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER60 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER60  (
    .ADR0(\BU2/U0/CHOICE3262 ),
    .ADR1(\BU2/U0/CHOICE3268 ),
    .ADR2(\BU2/U0/CHOICE3272 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0])
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER60/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .O(\BU2/U0/N66129 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker193971 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker193971  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_Ker193971/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/N66131 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194341 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194341  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194341/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/N66133 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194101 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194101  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194101/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .O(\BU2/U0/N66135 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78  (
    .ADR0(\BU2/U0/CHOICE2846 ),
    .ADR1(\BU2/U0/N65468 ),
    .ADR2(\BU2/U0/CHOICE2833 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_RESETb1/LUT2_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .O(\BU2/U0/N66138 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<4>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<0>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<1>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<2>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<3>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_TX_UNDERRUN_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER48/O ),
    .O(\BU2/U0/CHOICE3272 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [12]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [12]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<12>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [12])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [11]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<11>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [11])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [10]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<10>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [10])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<9>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [9])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<8>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<7>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<6>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005<5>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_271/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_27 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_261/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_26 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [13]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_231/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_23 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_241/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_24 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[3] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_251/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_25 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493_SW0/O ),
    .O(\BU2/U0/N51500 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR1(\BU2/U0/N66193 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05111/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0511 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR2(\BU2/U0/N66288 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04631/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0463 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0  (
    .ADR0(\BU2/U0/CHOICE2849 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>78_SW0/O ),
    .O(\BU2/U0/N65468 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04601/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0460 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0350 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04591/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0459 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04471/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0447 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0291 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04461/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0446 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_571/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_57 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_551/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_55 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_541/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_54 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_531/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_53 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032  (
    .ADR0(\BU2/U0/CHOICE2768 ),
    .ADR1(\BU2/U0/CHOICE2771 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035032/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0350 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TC_ASSIGN_I0 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_511/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_51 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_521/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_52 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_501/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_50 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65388 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141 .INIT = 16'hF800;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141  (
    .ADR0(\BU2/U0/CHOICE3126 ),
    .ADR1(\BU2/U0/CHOICE3129 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR3(\BU2/U0/CHOICE3132 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029141/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0291 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117  (
    .ADR0(\BU2/U0/N65873 ),
    .ADR1(\BU2/U0/CHOICE2870 ),
    .ADR2(\BU2/U0/CHOICE2881 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_END_OF_TX1 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_END_OF_TX1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR2(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_END_OF_TX )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_END_OF_TX1/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_END_OF_TX ),
    .O(\BU2/U0/N66180 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_561/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_56 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[14] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[5] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<5>16_SW0/O ),
    .O(\BU2/U0/N65388 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DELAYED ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0179 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01731 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01731  (
    .ADR0(\BU2/U0/N66216 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0173 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01731/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0173 ),
    .O(\BU2/U0/N66185 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL1 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL1/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL ),
    .O(\BU2/U0/N66187 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [10]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194041 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194041  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194041/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .O(\BU2/U0/N66190 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [12]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID1 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0273 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID1/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID ),
    .O(\BU2/U0/N66193 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING1 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING1/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .O(\BU2/U0/N66195 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [1]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4470 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [2]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4474 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [3]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4478 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [4]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4482 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [5]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4486 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [6]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4490 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [7]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4494 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [8]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4498 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [9]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4502 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [10]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4506 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [11]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4510 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [12]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4514 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [13]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4518 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4542 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [2]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4548 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4562 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>lut/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4566 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [14]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215181 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215181  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21520 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215181/LUT3_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21520 ),
    .O(\BU2/U0/N66216 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [11]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221 .INIT = 16'h3B08;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/N66102 ),
    .ADR2(tieemacconfigvec_7[65]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_221/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_22 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt_11 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt_11  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021 .INIT = 16'h000E;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker229021/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22904 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00071 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00071  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00071/LUT2_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .O(\BU2/U0/N66231 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209 .INIT = 16'hFF27;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY [2]),
    .ADR2(\BU2/U0/N65527 ),
    .ADR3(\BU2/U0/CHOICE3208 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1 .INIT = 16'hAEA2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02564/O ),
    .O(\BU2/U0/CHOICE3115 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_271/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_27 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221 .INIT = 16'h3B08;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/N66312 ),
    .ADR2(tieemacconfigvec_7[65]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_221/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_22 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_231/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_23 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[3] ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_251/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_25 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65392 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[13] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[4] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<4>16_SW0/O ),
    .O(\BU2/U0/N65392 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50/O ),
    .O(\BU2/U0/CHOICE1830 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324_12 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324_12  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ),
    .ADR3(\BU2/U0/N53310 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324 ),
    .O(\BU2/U0/N66248 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00921 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00921  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0092 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00921/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0092 ),
    .O(\BU2/U0/N66250 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161261/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16128 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01021 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01021  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0102 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01021/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0102 ),
    .O(\BU2/U0/N66253 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01011 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01011  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01011/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ),
    .O(\BU2/U0/N66255 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841  (
    .ADR0(\BU2/U0/N66255 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00841/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0084 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00821/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0082 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00811/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0081 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00801/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0080 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00791/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0079 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00781/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0078 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .ADR3(\BU2/U0/N66253 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00861/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0086 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0102 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00701/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0070 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/N66250 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00611/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0061 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16128 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00601/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0060 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00581/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0058 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00571/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0057 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0092 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00561/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0056 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0092 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00471/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0047 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00461/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0046 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0101 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00451/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0045 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_581/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_58 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR1(\BU2/U0/CHOICE3136 ),
    .ADR2(\BU2/U0/CHOICE3141 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046140/O ),
    .O(\BU2/U0/CHOICE3145 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt_13 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt_13  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [0]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n00001/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00771/O ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0077 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65396 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[12] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[3] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<3>16_SW0/O ),
    .O(\BU2/U0/N65396 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1_14 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1_14  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [4]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt_15 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt_15  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [3]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN_SW0/O ),
    .O(\BU2/U0/N53520 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1_16 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1_16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [5]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O ),
    .O(\BU2/U0/CHOICE1790 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_SW0/O ),
    .O(\BU2/U0/N53474 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65400 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[11] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[2] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<2>16_SW0/O ),
    .O(\BU2/U0/N65400 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197_17 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197_17  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .ADR3(\BU2/U0/N53310 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197 ),
    .O(\BU2/U0/N66288 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_18 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS_18  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .ADR3(\BU2/U0/N53474 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ),
    .O(\BU2/U0/N66290 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I259  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C4 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I259/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I259/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I259/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C5 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I272  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C5 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I272/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I272/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I272/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I285  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C6 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I285/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I285/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I285/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I246  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C3 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I246/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I246/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I246/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I233  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C2 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I233/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I233/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I233/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I26  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I26/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I26/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I26/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I4  (
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I4/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I4/MUXCY_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I4/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TC_ASSIGN_I0 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt_19 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt_19  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [2]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071_SW0/O ),
    .O(\BU2/U0/N52594 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21 .INIT = 8'h90;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE1819 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21/O ),
    .O(\BU2/U0/CHOICE1820 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN .INIT = 16'h5554;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE [0]),
    .ADR3(\BU2/U0/N53520 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0])
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EN/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .O(\BU2/U0/N66295 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0068_20 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0068_20  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX__n0046 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR2(\BU2/U0/N53563 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0068 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0068/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0068 ),
    .O(\BU2/U0/N66297 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt_21 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt_21  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [4]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65404 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[10] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[1] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<1>16_SW0/O ),
    .O(\BU2/U0/N65404 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1_22 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1_22  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [3]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65280 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16092 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087_SW0/O ),
    .O(\BU2/U0/N51803 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[16] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[7] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<7>16_SW0/O ),
    .O(\BU2/U0/N65280 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199 .INIT = 16'h00AE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199  (
    .ADR0(\BU2/U0/CHOICE1791 ),
    .ADR1(\BU2/U0/CHOICE1804 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O ),
    .O(\BU2/U0/CHOICE1809 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109/O ),
    .O(\BU2/U0/CHOICE1844 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199 .INIT = 16'h00AE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199  (
    .ADR0(\BU2/U0/CHOICE1685 ),
    .ADR1(\BU2/U0/CHOICE1698 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>199/O ),
    .O(\BU2/U0/CHOICE1703 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>117/O ),
    .O(\BU2/U0/CHOICE1684 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N65284 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<6>16/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt_23 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt_23  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [6]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN__n0005 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN__n0005  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [0]),
    .ADR3(\BU2/U0/N65067 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN__n0005/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .O(\BU2/U0/N66312 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84  (
    .ADR0(\BU2/U0/CHOICE3082 ),
    .ADR1(\BU2/U0/N65368 ),
    .ADR2(\BU2/U0/CHOICE3085 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149  (
    .ADR0(\BU2/U0/CHOICE2720 ),
    .ADR1(\BU2/U0/CHOICE2752 ),
    .ADR2(\BU2/U0/CHOICE2726 ),
    .ADR3(\BU2/U0/N65350 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296_24 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296_24  (
    .ADR0(\BU2/U0/N61770 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker214981 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker214981  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker214981/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .O(\BU2/U0/N66317 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/CHOICE3067 ),
    .ADR2(\BU2/U0/CHOICE3073 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>84_SW0/O ),
    .O(\BU2/U0/N65368 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354_25 .INIT = 16'hAAEF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354_25  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR2(\BU2/U0/N62536 ),
    .ADR3(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84  (
    .ADR0(\BU2/U0/CHOICE3106 ),
    .ADR1(\BU2/U0/N65372 ),
    .ADR2(\BU2/U0/CHOICE3109 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/CHOICE3091 ),
    .ADR2(\BU2/U0/CHOICE3097 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>84_SW0/O ),
    .O(\BU2/U0/N65372 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77  (
    .ADR0(\BU2/U0/CHOICE3058 ),
    .ADR1(\BU2/U0/N65376 ),
    .ADR2(\BU2/U0/CHOICE3061 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER11/O ),
    .O(\BU2/U0/CHOICE3259 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0  (
    .ADR0(\BU2/U0/CHOICE2735 ),
    .ADR1(\BU2/U0/CHOICE2730 ),
    .ADR2(\BU2/U0/CHOICE2716 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>149_SW0/O ),
    .O(\BU2/U0/N65350 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/CHOICE3044 ),
    .ADR2(\BU2/U0/CHOICE3050 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>77_SW0/O ),
    .O(\BU2/U0/N65376 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>21/O ),
    .O(\BU2/U0/CHOICE2839 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1_26 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1_26  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [6]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58_SW0/O ),
    .O(\BU2/U0/N65743 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000057 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000057  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [0]),
    .ADR1(\BU2/U0/N65878 ),
    .ADR2(\BU2/U0/CHOICE2673 ),
    .ADR3(\BU2/U0/CHOICE2680 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000057/LUT4_D_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 ),
    .O(\BU2/U0/N66330 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [14]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58_SW0/O ),
    .O(\BU2/U0/N65747 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_TX_END_OF_TX ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16_SW0/O ),
    .O(\BU2/U0/N65424 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212  (
    .ADR0(\BU2/U0/CHOICE2899 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046212/O ),
    .O(\BU2/U0/CHOICE2900 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28  (
    .ADR0(\BU2/U0/CHOICE2987 ),
    .ADR1(\BU2/U0/CHOICE2994 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28/LUT2_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In28/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1  (
    .ADR0(\BU2/U0/CHOICE2863 ),
    .ADR1(\BU2/U0/CHOICE2867 ),
    .ADR2(\BU2/U0/CHOICE2857 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>117_SW1/O ),
    .O(\BU2/U0/N65873 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77  (
    .ADR0(\BU2/U0/CHOICE3012 ),
    .ADR1(\BU2/U0/N65380 ),
    .ADR2(\BU2/U0/CHOICE3015 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT ),
    .ADR2(\BU2/U0/N65424 ),
    .ADR3(\BU2/U0/CHOICE2688 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In16/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n004610 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n004610  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX__n0067 ),
    .ADR3(\BU2/U0/CHOICE1379 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n004610/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n004610/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n004610/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0046 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022__n0002 ),
    .ADR2(\BU2/U0/CHOICE3237 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0/LUT3_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010209_SW0/O ),
    .O(\BU2/U0/N65527 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt_27 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt_27  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [5]),
    .ADR1(GND),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt/LUT1_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt/O ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77  (
    .ADR0(\BU2/U0/CHOICE3035 ),
    .ADR1(\BU2/U0/N65384 ),
    .ADR2(\BU2/U0/CHOICE3038 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77/O ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/CHOICE2998 ),
    .ADR2(\BU2/U0/CHOICE3004 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>77_SW0/O ),
    .O(\BU2/U0/N65380 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/CHOICE3021 ),
    .ADR2(\BU2/U0/CHOICE3027 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>77_SW0/O ),
    .O(\BU2/U0/N65384 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9 .INIT = 16'hF200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX__n0067 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_CONTROL_COMPLETE ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In9/O ),
    .O(\BU2/U0/CHOICE2987 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX__n0067 ),
    .ADR3(\BU2/U0/CHOICE1379 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1/O )
  );
  X_BUF \BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1/LUT4_L_BUF  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n004610_1/O ),
    .O(\BU2/U0/N66008 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>67_F .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>67_F  (
    .ADR0(\BU2/U0/CHOICE2875 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19418 ),
    .O(\BU2/U0/N66097 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>67  (
    .IA(\BU2/U0/N66097 ),
    .IB(\BU2/U0/N66099 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .O(\BU2/U0/CHOICE2881 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<10>161_F .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<10>161_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [1]),
    .O(\BU2/U0/N66092 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<10>161  (
    .IA(\BU2/U0/N66092 ),
    .IB(\BU2/U0/N66094 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [10]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [10])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010212_F .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010212_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR1(\BU2/U0/CHOICE3286 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY [1]),
    .ADR3(\BU2/U0/CHOICE3315 ),
    .O(\BU2/U0/N66087 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010212  (
    .IA(\BU2/U0/N66087 ),
    .IB(\BU2/U0/N66089 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<11>161_F .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<11>161_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [2]),
    .O(\BU2/U0/N66082 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<11>161  (
    .IA(\BU2/U0/N66082 ),
    .IB(\BU2/U0/N66084 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [11]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [11])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>161_F .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>161_F  (
    .ADR0(\BU2/U0/CHOICE1945 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [3]),
    .O(\BU2/U0/N66077 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>161  (
    .IA(\BU2/U0/N66077 ),
    .IB(\BU2/U0/N66079 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [9])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_FORCE_QUIET_Result16_F .INIT = 16'h000E;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_FORCE_QUIET_Result16_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .O(\BU2/U0/N66072 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_FORCE_QUIET_Result16  (
    .IA(\BU2/U0/N66072 ),
    .IB(\BU2/U0/N66074 ),
    .SEL(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<12>161_F .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<12>161_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [3]),
    .O(\BU2/U0/N66067 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<12>161  (
    .IA(\BU2/U0/N66067 ),
    .IB(\BU2/U0/N66069 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [12]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [12])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<14>161_F .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<14>161_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [5]),
    .O(\BU2/U0/N66062 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<14>161  (
    .IA(\BU2/U0/N66062 ),
    .IB(\BU2/U0/N66064 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [14]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [14])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<13>161_F .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<13>161_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [4]),
    .O(\BU2/U0/N66057 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<13>161  (
    .IA(\BU2/U0/N66057 ),
    .IB(\BU2/U0/N66059 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [13]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [13])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_F .INIT = 16'h1D45;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/N66052 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80  (
    .IA(\BU2/U0/N66052 ),
    .IB(\BU2/U0/N66054 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .O(\BU2/U0/CHOICE1677 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result43_F .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result43_F  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxer),
    .ADR2(\BU2/U0/CHOICE2628 ),
    .O(\BU2/U0/N66047 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result43  (
    .IA(\BU2/U0/N66047 ),
    .IB(\BU2/U0/N66049 ),
    .SEL(\BU2/U0/CHOICE2633 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RX_ER )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_F .INIT = 16'h1D45;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/N66042 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80  (
    .IA(\BU2/U0/N66042 ),
    .IB(\BU2/U0/N66044 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .O(\BU2/U0/CHOICE1783 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_F .INIT = 16'h0006;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/N66037 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192  (
    .IA(\BU2/U0/N66037 ),
    .IB(\BU2/U0/N66039 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/CHOICE1863 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_Mmux__n0029_Result34_F .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_Mmux__n0029_Result34_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/N66032 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_Mmux__n0029_Result34  (
    .IA(\BU2/U0/N66032 ),
    .IB(\BU2/U0/N66034 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0029 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_F .INIT = 16'h0006;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_F  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/N66027 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192  (
    .IA(\BU2/U0/N66027 ),
    .IB(\BU2/U0/N66029 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/CHOICE1757 )
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7_28 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7_28  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9_29 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9_29  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8_30 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8_30  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7_31 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7_31  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6_32 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6_32  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5_33 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5_33  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4_34 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4_34  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3_35 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3_35  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2_36 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2_36  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1_37 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1_37  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 )
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6_38 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6_38  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5_39 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5_39  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4_40 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4_40  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3_41 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3_41  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2_42 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2_42  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1_43 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1_43  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1_44 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1_44  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1_45 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1_45  (
    .I(\BU2/U0/N66008 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0068 ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1_46 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1_46  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0076 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0462 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1_47 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1_47  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0443 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1_48 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1_48  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt_49 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt_49  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt_50 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt_50  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt_51 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt_51  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt_52 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt_52  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt_53 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt_53  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt_54 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt_54  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt_55 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt_55  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt_56 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt_56  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt_57 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt_57  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010116 .INIT = 16'h0281;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010116  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/CHOICE3232 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148856 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148856  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [5]),
    .ADR1(\BU2/U0/N65882 ),
    .ADR2(\BU2/U0/CHOICE2974 ),
    .ADR3(\BU2/U0/CHOICE2981 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21490 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [17]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [25]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/CHOICE3073 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>55 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>55  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [35]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [43]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .O(\BU2/U0/CHOICE2849 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt_58 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt_58  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001023 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001023  (
    .ADR0(\BU2/U0/CHOICE3280 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [5]),
    .ADR3(\BU2/U0/N65436 ),
    .O(\BU2/U0/CHOICE3286 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010150_SW0 .INIT = 16'hE7FF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010150_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/N65487 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>30 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>30  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [23]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .O(\BU2/U0/CHOICE2867 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt_59 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt_59  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00120 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX__n00120  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/CHOICE2590 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [22]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [30]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/CHOICE3097 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG38 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG38  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .ADR1(\BU2/U0/N65432 ),
    .ADR2(\BU2/U0/CHOICE2587 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In9 .INIT = 16'hA2AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In9  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/CHOICE2688 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>15  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [3]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2804 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In21_SW0 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In21_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .O(\BU2/U0/N65416 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt_60 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt_60  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029114 .INIT = 16'h0DFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029114  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .O(\BU2/U0/CHOICE3126 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012144 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012144  (
    .ADR0(\BU2/U0/N65464 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE3161 ),
    .ADR3(\BU2/U0/CHOICE3182 ),
    .O(\BU2/U0/CHOICE3193 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG28 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG28  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [3]),
    .O(\BU2/U0/CHOICE2587 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In21 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR2(\BU2/U0/N65416 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/CHOICE2994 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [21]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [29]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/CHOICE3027 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010150 .INIT = 16'h7F5D;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010150  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22745 ),
    .ADR2(\BU2/U0/N65487 ),
    .ADR3(\BU2/U0/CHOICE3232 ),
    .O(\BU2/U0/CHOICE3237 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>15  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [0]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2826 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_G .INIT = 16'h0070;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/N66029 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>61 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>61  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [16]),
    .O(\BU2/U0/CHOICE2735 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00085 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00085  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH ),
    .O(\BU2/U0/CHOICE2693 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>40 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>40  (
    .ADR0(\BU2/U0/CHOICE2839 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .ADR2(\BU2/U0/CHOICE2844 ),
    .O(\BU2/U0/CHOICE2846 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt_61 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt_61  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012144 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012144  (
    .ADR0(\BU2/U0/N65460 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE2908 ),
    .ADR3(\BU2/U0/CHOICE2929 ),
    .O(\BU2/U0/CHOICE2940 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt_62 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt_62  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035012 .INIT = 8'h8F;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n035012  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ),
    .ADR2(\BU2/U0/N66195 ),
    .O(\BU2/U0/CHOICE2771 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001218 .INIT = 8'h06;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001218  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/CHOICE3161 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465_63 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465_63  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR1(\BU2/U0/N61129 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG38_SW0 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG38_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [6]),
    .O(\BU2/U0/N65432 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465_SW0 .INIT = 16'hFBBB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .O(\BU2/U0/N61129 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt_64 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt_64  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021834_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021834_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [8]),
    .O(\BU2/U0/N65428 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt_65 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt_65  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt_66 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt_66  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt_67 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt_67  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [15]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [7]),
    .ADR3(\BU2/U0/N66133 ),
    .O(\BU2/U0/CHOICE2863 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>32 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>32  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [27]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [19]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/CHOICE2844 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>57 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>57  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [12]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/CHOICE3058 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01441 .INIT = 16'h0BBB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01441  (
    .ADR0(\BU2/U0/N53281 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0144 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>50 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>50  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [32]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .O(\BU2/U0/CHOICE2730 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03507 .INIT = 8'h23;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03507  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .O(\BU2/U0/CHOICE2768 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt_68 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt_68  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04451 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04451  (
    .ADR0(\BU2/U0/CHOICE2785 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR3(\BU2/U0/CHOICE2778 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0445 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<3>0  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [3]),
    .O(\BU2/U0/CHOICE2798 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001218 .INIT = 8'h06;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001218  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/CHOICE2908 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046216 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046216  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0177 ),
    .ADR1(\BU2/U0/CHOICE2900 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0462 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00455 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00455  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [3]),
    .O(\BU2/U0/CHOICE3246 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047583 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047583  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/CHOICE2553 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL ),
    .ADR3(\BU2/U0/N65440 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0475 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt_69 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt_69  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [36]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [44]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .O(\BU2/U0/CHOICE3044 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result12 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result12  (
    .ADR0(\BU2/U0/CHOICE2632 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .O(\BU2/U0/CHOICE2633 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<0>0  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [0]),
    .O(\BU2/U0/CHOICE2820 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt_70 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt_70  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>62 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>62  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [12]),
    .O(\BU2/U0/CHOICE3061 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt_71 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt_71  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result8 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result8  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3 ),
    .O(\BU2/U0/CHOICE2632 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001015 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001015  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [7]),
    .O(\BU2/U0/CHOICE3205 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n004511 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n004511  (
    .ADR0(\BU2/U0/CHOICE3246 ),
    .ADR1(\BU2/U0/CHOICE3205 ),
    .O(\BU2/U0/CHOICE3250 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>40 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>40  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/CHOICE2726 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04614 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04614  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ),
    .O(\BU2/U0/CHOICE3136 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>58  (
    .ADR0(\BU2/U0/N65747 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .O(\BU2/U0/CHOICE3106 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt_72 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt_72  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt_73 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt_73  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1 ),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2628 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000045 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000045  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [8]),
    .O(\BU2/U0/CHOICE2680 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt_74 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt_74  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n001223 .INIT = 8'h57;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n001223  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT ),
    .O(\BU2/U0/CHOICE2600 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>58  (
    .ADR0(\BU2/U0/N65743 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .O(\BU2/U0/CHOICE3082 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt_75 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt_75  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1_76 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1_76  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt_77 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt_77  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010107 .INIT = 16'h0281;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010107  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/CHOICE3310 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148844 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148844  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [14]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [13]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [1]),
    .O(\BU2/U0/CHOICE2981 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04629 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04629  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR2(\BU2/U0/N66187 ),
    .O(\BU2/U0/CHOICE2899 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001033 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001033  (
    .ADR0(\BU2/U0/CHOICE3246 ),
    .ADR1(\BU2/U0/CHOICE3205 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .O(\BU2/U0/CHOICE3208 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010141_SW0 .INIT = 16'hE7FF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010141_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .O(\BU2/U0/N65483 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>15  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [2]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2793 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [37]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [45]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .O(\BU2/U0/CHOICE3021 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047532 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047532  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [1]),
    .O(\BU2/U0/CHOICE2560 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001248 .INIT = 16'h9D80;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001248  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/CHOICE3171 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>68 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>68  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [14]),
    .O(\BU2/U0/CHOICE3109 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012144_SW0 .INIT = 16'hFF06;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012144_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22745 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .ADR3(\BU2/U0/CHOICE3171 ),
    .O(\BU2/U0/N65464 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148831 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148831  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [12]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [15]),
    .O(\BU2/U0/CHOICE2974 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001290 .INIT = 16'hFF90;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001290  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/CHOICE2928 ),
    .O(\BU2/U0/CHOICE2929 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046115 .INIT = 16'h000E;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046115  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .O(\BU2/U0/CHOICE3141 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>18 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>18  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [40]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .O(\BU2/U0/CHOICE2720 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>68 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>68  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [9]),
    .O(\BU2/U0/CHOICE3085 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010141 .INIT = 16'h7F5D;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010141  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22745 ),
    .ADR2(\BU2/U0/N65483 ),
    .ADR3(\BU2/U0/CHOICE3310 ),
    .O(\BU2/U0/CHOICE3315 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000032 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000032  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [4]),
    .O(\BU2/U0/CHOICE2673 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt_78 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt_78  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt_79 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt_79  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>52 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>52  (
    .ADR0(\BU2/U0/N66131 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [31]),
    .O(\BU2/U0/CHOICE2875 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt_80 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt_80  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [18]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [26]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/CHOICE3004 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>15  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [1]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2815 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047583_SW0 .INIT = 16'h1800;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047583_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [9]),
    .ADR3(\BU2/U0/CHOICE2560 ),
    .O(\BU2/U0/N65440 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_Mmux__n0029_Result34_G .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_Mmux__n0029_Result34_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_IFG_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .O(\BU2/U0/N66034 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047513 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n047513  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [8]),
    .O(\BU2/U0/CHOICE2553 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00011 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER21 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER21  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR1(\BU2/U0/CHOICE3259 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION ),
    .O(\BU2/U0/CHOICE3262 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [15]),
    .O(\BU2/U0/CHOICE2857 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_321 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_321  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_32 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296_SW0 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ),
    .O(\BU2/U0/N61770 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354_SW0 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .O(\BU2/U0/N62536 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<2>0  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [2]),
    .O(\BU2/U0/CHOICE2787 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt_81 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt_81  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt_82 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt_82  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN__n0005_SW0 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN__n0005_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [4]),
    .O(\BU2/U0/N65067 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt_83 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt_83  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021834 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021834  (
    .ADR0(\BU2/U0/CHOICE2949 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [1]),
    .ADR3(\BU2/U0/N65428 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0218 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n028726 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n028726  (
    .ADR0(\BU2/U0/CHOICE2778 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR2(\BU2/U0/CHOICE2785 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0287 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001175_SW0 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001175_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [9]),
    .O(\BU2/U0/N65358 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In25 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In25  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ),
    .O(\BU2/U0/CHOICE2389 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [1]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65500 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000962 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000962  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD ),
    .O(\BU2/U0/CHOICE2409 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In46_SW0 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In46_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 ),
    .O(\BU2/U0/N65472 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003321 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003321  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [6]),
    .O(\BU2/U0/CHOICE2117 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001175 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001175  (
    .ADR0(\BU2/U0/CHOICE2494 ),
    .ADR1(\BU2/U0/CHOICE2501 ),
    .ADR2(\BU2/U0/CHOICE2486 ),
    .ADR3(\BU2/U0/N65358 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0011 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001223 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001223  (
    .ADR0(\BU2/U0/CHOICE2080 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>30 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>30  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/CHOICE2152 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In32 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In32  (
    .ADR0(\BU2/U0/N65448 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_N21825 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2 ),
    .ADR3(\BU2/U0/CHOICE2157 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01716 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01716  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ),
    .O(\BU2/U0/CHOICE2436 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00149 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00149  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [13]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [15]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [1]),
    .O(\BU2/U0/CHOICE2041 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336_SW0 .INIT = 16'hFBBB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/N59896 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001216 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001216  (
    .ADR0(\BU2/U0/CHOICE2079 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .O(\BU2/U0/CHOICE2080 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336_84 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336_84  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_COL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR3(\BU2/U0/N59896 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker168977 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker168977  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [1]),
    .O(\BU2/U0/CHOICE2257 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [2]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2373 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG62 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG62  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [16]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [17]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [18]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/CHOICE2250 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001212 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n001212  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ),
    .O(\BU2/U0/CHOICE2079 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00144 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00144  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [10]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [11]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [12]),
    .O(\BU2/U0/CHOICE2038 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt_85 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt_85  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n016121 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n016121  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN ),
    .ADR1(\BU2/U0/N65444 ),
    .ADR2(\BU2/U0/CHOICE2277 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010415 .INIT = 16'h007F;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010415  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .O(\BU2/U0/CHOICE2185 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE57 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE57  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [9]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [14]),
    .O(\BU2/U0/CHOICE2470 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG17 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG17  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [9]),
    .ADR3(\BU2/U0/N65412 ),
    .O(\BU2/U0/CHOICE2230 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE69_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE69_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [13]),
    .O(\BU2/U0/N65330 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt_86 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt_86  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt_87 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt_87  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n012810 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n012810  (
    .ADR0(\BU2/U0/CHOICE2031 ),
    .ADR1(\BU2/U0/CHOICE2034 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0128 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001127 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001127  (
    .ADR0(\BU2/U0/CHOICE2211 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [0]),
    .O(\BU2/U0/CHOICE2216 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01289 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01289  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7 ),
    .O(\BU2/U0/CHOICE2034 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005118 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005118  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16087 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH ),
    .O(\BU2/U0/CHOICE2201 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003331_SW0 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003331_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [7]),
    .O(\BU2/U0/N65452 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE69 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE69  (
    .ADR0(\BU2/U0/CHOICE2455 ),
    .ADR1(\BU2/U0/CHOICE2463 ),
    .ADR2(\BU2/U0/CHOICE2470 ),
    .ADR3(\BU2/U0/N65330 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt_88 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt_88  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt_89 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt_89  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [2]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2313 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n017117 .INIT = 16'h22F2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n017117  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .O(\BU2/U0/CHOICE2441 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01284 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01284  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3 ),
    .O(\BU2/U0/CHOICE2031 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt_90 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt_90  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>43 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>43  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [47]),
    .O(\BU2/U0/CHOICE2870 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [3]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2337 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [0]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2361 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In16 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .O(\BU2/U0/CHOICE2162 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00092 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00092  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [10]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16530 ),
    .O(\BU2/U0/CHOICE2394 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker1689718 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker1689718  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [2]),
    .O(\BU2/U0/CHOICE2262 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [0]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65496 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013010 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013010  (
    .ADR0(\BU2/U0/CHOICE2024 ),
    .ADR1(\BU2/U0/CHOICE2027 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0130 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n017125 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n017125  (
    .ADR0(\BU2/U0/CHOICE2436 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR2(\BU2/U0/CHOICE2441 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0171 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01309 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01309  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7 ),
    .O(\BU2/U0/CHOICE2027 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_DV_Result16 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_DV_Result16  (
    .ADR0(\BU2/U0/CHOICE1120 ),
    .ADR1(corehassgmii),
    .ADR2(phyemacrxdv),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RX_DV )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n002124 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n002124  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_DATA [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_DATA [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_DATA [7]),
    .O(\BU2/U0/CHOICE2516 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [1]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2349 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt_91 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt_91  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003430 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003430  (
    .ADR0(\BU2/U0/CHOICE2104 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [1]),
    .ADR3(\BU2/U0/N65456 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0034 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In_92 .INIT = 16'hF800;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In_92  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ),
    .ADR1(\BU2/U0/N58329 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_N21825 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In_SW0 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .O(\BU2/U0/N58329 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01304 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01304  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3 ),
    .O(\BU2/U0/CHOICE2024 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [0]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2301 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG37 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG37  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [10]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [11]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [12]),
    .O(\BU2/U0/CHOICE2237 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt_93 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt_93  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00518 .INIT = 8'h07;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00518  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE ),
    .O(\BU2/U0/CHOICE2197 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt_94 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt_94  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt_95 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt_95  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003420 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003420  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [6]),
    .O(\BU2/U0/CHOICE2104 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [3]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2289 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n012910 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n012910  (
    .ADR0(\BU2/U0/CHOICE2017 ),
    .ADR1(\BU2/U0/CHOICE2020 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0129 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt_96 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt_96  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01299 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01299  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .O(\BU2/U0/CHOICE2020 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In32_SW0 .INIT = 8'hBF;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In32_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR1(\BU2/U0/CHOICE2162 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ),
    .O(\BU2/U0/N65448 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [3]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65508 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In4 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In4  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .O(\BU2/U0/CHOICE2157 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01619 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01619  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [7]),
    .O(\BU2/U0/CHOICE2277 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001114 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001114  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [1]),
    .O(\BU2/U0/CHOICE2211 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt_97 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt_97  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In27 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In27  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT ),
    .O(\BU2/U0/CHOICE2177 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01294 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01294  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .O(\BU2/U0/CHOICE2017 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n016121_SW0 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n016121_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [3]),
    .O(\BU2/U0/N65444 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [7]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65492 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012144_SW0 .INIT = 16'hFF06;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012144_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22745 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .ADR3(\BU2/U0/CHOICE2918 ),
    .O(\BU2/U0/N65460 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n002148 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n002148  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [3]),
    .O(\BU2/U0/CHOICE2524 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n025614 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n025614  (
    .ADR0(\BU2/U0/CHOICE3115 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [2]),
    .ADR3(\BU2/U0/N65420 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03194 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03194  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .O(\BU2/U0/CHOICE2424 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059_98 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059_98  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16092 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR3(\BU2/U0/N57931 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059_SW0 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [1]),
    .O(\BU2/U0/N57931 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013110 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013110  (
    .ADR0(\BU2/U0/CHOICE2010 ),
    .ADR1(\BU2/U0/CHOICE2013 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0131 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04661 .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04661  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0218 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01319 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01319  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7 ),
    .O(\BU2/U0/CHOICE2013 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001125 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001125  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [11]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [12]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [13]),
    .O(\BU2/U0/CHOICE2486 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [6]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65520 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001111 .INIT = 16'hFF7F;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001111  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [3]),
    .O(\BU2/U0/CHOICE2209 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003430_SW0 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003430_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [3]),
    .O(\BU2/U0/N65456 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0015_99 .INIT = 16'h7776;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0015_99  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/N65764 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0015 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0015_SW1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0015_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .O(\BU2/U0/N65764 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n002022 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n002022  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/CHOICE2122 ),
    .ADR2(\BU2/U0/CHOICE2126 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01314 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01314  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3 ),
    .O(\BU2/U0/CHOICE2010 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt_100 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt_100  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010435 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010435  (
    .ADR0(\BU2/U0/CHOICE2191 ),
    .ADR1(\BU2/U0/CHOICE2185 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0104 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>22 .INIT = 16'hF078;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>22  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [4]),
    .ADR3(\BU2/U0/N65751 ),
    .O(\BU2/U0/CHOICE2152 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt_101 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt_101  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE21 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE21  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [3]),
    .O(\BU2/U0/CHOICE2455 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [2]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65504 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In13 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In13  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .ADR3(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .O(\BU2/U0/CHOICE2384 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n002161 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n002161  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [7]),
    .O(\BU2/U0/CHOICE2531 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013210 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n013210  (
    .ADR0(\BU2/U0/CHOICE2003 ),
    .ADR1(\BU2/U0/CHOICE2006 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0132 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000921 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000921  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .O(\BU2/U0/CHOICE2403 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01329 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01329  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7 ),
    .O(\BU2/U0/CHOICE2006 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n002174_SW0 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n002174_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_DATA [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_DATA [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_DATA [0]),
    .O(\BU2/U0/N65354 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n002012 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n002012  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .O(\BU2/U0/CHOICE2126 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG17_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG17_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [13]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [15]),
    .O(\BU2/U0/N65412 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt_102 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt_102  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013<1>0  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [1]),
    .O(\BU2/U0/CHOICE2809 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010432 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n010432  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256 ),
    .O(\BU2/U0/CHOICE2191 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n002174 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n002174  (
    .ADR0(\BU2/U0/CHOICE2524 ),
    .ADR1(\BU2/U0/CHOICE2531 ),
    .ADR2(\BU2/U0/CHOICE2516 ),
    .ADR3(\BU2/U0/N65354 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0021 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01324 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01324  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3 ),
    .O(\BU2/U0/CHOICE2003 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005419 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005419  (
    .ADR0(\BU2/U0/CHOICE2085 ),
    .ADR1(\BU2/U0/CHOICE2091 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0054 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In11 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In11  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .O(\BU2/U0/CHOICE2173 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005416 .INIT = 16'hFBBB;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005416  (
    .ADR0(\BU2/U0/CHOICE2087 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .O(\BU2/U0/CHOICE2091 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>57 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>57  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [13]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/CHOICE3035 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>22_SW0 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<4>22_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .O(\BU2/U0/N65751 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001149 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001149  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [14]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [15]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17 ),
    .O(\BU2/U0/CHOICE2494 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n031914 .INIT = 16'h0888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n031914  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .O(\BU2/U0/CHOICE2430 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2> .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/N50904 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004_103 .INIT = 16'hDCD0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004_103  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .ADR3(\BU2/U0/N50382 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004_SW0 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1 ),
    .O(\BU2/U0/N50382 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>_SW0 .INIT = 8'h95;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [0]),
    .O(\BU2/U0/N50904 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_G .INIT = 16'h0070;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>192_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/N66039 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0058_Result_SW1 .INIT = 8'h96;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0058_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .O(\BU2/U0/N65788 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458_104 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458_104  (
    .ADR0(\BU2/U0/N52476 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21520 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>59 .INIT = 16'h1800;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>59  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .ADR3(\BU2/U0/CHOICE1724 ),
    .O(\BU2/U0/CHOICE1725 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458_SW0 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0174 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ),
    .O(\BU2/U0/N52476 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0060_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0060_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0296 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .O(\BU2/U0/N65792 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>213 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>213  (
    .ADR0(\BU2/U0/CHOICE1703 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE1677 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0060_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0060_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0297 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65792 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0060 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>120 .INIT = 16'h9200;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>120  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .ADR3(\BU2/U0/CHOICE1844 ),
    .O(\BU2/U0/CHOICE1845 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0062_Result_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0062_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .O(\BU2/U0/N65946 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015_105 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015_105  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/N65808 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024_106 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024_106  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16530 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .ADR3(\BU2/U0/N50348 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .O(\BU2/U0/N50348 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015_SW1 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ),
    .O(\BU2/U0/N65808 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0087  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/N51803 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_BYTE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>213 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>213  (
    .ADR0(\BU2/U0/CHOICE1809 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE1783 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt_107 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt_107  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>122 .INIT = 16'h8B00;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>122  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/CHOICE1684 ),
    .O(\BU2/U0/CHOICE1685 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_G .INIT = 16'h1D3C;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/N66044 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt_108 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt_108  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029138 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029138  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE ),
    .O(\BU2/U0/CHOICE3132 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0062_Result .INIT = 16'h2EE2;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0062_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0299 [1]),
    .ADR3(\BU2/U0/N65946 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0062 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_DV_Result15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_DV_Result15  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3 ),
    .ADR3(corehassgmii),
    .O(\BU2/U0/CHOICE1120 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<3> .INIT = 16'h2772;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<3>  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [3]),
    .ADR3(\BU2/U0/N52276 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017_109 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017_109  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .ADR2(\BU2/U0/N50321 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017_SW0 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .O(\BU2/U0/N50321 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2> .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/N51126 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>_SW0 .INIT = 8'h95;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [0]),
    .O(\BU2/U0/N51126 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt_110 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt_110  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<3>_SW0 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<3>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [1]),
    .O(\BU2/U0/N52276 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0062_Result .INIT = 16'h2EE2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0062_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0299 [1]),
    .ADR3(\BU2/U0/N65942 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0062 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0062_Result_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0062_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .O(\BU2/U0/N65942 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0063_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0063_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0299 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .O(\BU2/U0/N65636 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt_111 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt_111  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<3> .INIT = 16'h00A9;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<3>  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .ADR1(\BU2/U0/N51423 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<3>_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<3>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .O(\BU2/U0/N51423 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0063_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0063_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65636 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0063 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt_112 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt_112  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0058_Result .INIT = 16'h2EE2;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0058_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 [1]),
    .ADR3(\BU2/U0/N65788 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0058 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016_113 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016_113  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .ADR2(\BU2/U0/N50294 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016_SW0 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ),
    .O(\BU2/U0/N50294 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0060_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0060_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0297 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0296 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .O(\BU2/U0/N65784 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0061_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0061_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65965 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0061 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<9>_rt_114 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<9>_rt_114  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<9>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt_115 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt_115  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt_116 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt_116  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0064_Result .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0064_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/N65961 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0064 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In_117 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In_117  (
    .ADR0(\BU2/U0/N50272 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS ),
    .ADR1(tieemacconfigvec_7[55]),
    .O(\BU2/U0/N50272 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014_118 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014_118  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ),
    .ADR3(\BU2/U0/N50821 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00661 .INIT = 16'hFF7F;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n00661  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR2(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0066 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0064_Result_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0064_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .O(\BU2/U0/N65961 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt_119 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt_119  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0064_Result .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0064_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR1(\BU2/U0/N65957 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0064 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0064_Result_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0064_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .O(\BU2/U0/N65957 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>16 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/CHOICE1819 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt_120 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt_120  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>21 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<4>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [20]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [28]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19399 ),
    .O(\BU2/U0/CHOICE3050 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0037 .INIT = 16'h222A;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0037  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .ADR3(\BU2/U0/N52831 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0037_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0037_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/N52831 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker16071  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR3(\BU2/U0/N52594 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt_121 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt_121  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt_122 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt_122  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt_123 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt_123  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt_124 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt_124  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<2> .INIT = 16'h8DD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [2]),
    .ADR3(\BU2/U0/N51935 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<2>_SW0 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .O(\BU2/U0/N51935 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190_125 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190_125  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR3(\BU2/U0/N50226 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/N50226 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt_126 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt_126  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014_127 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014_127  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .ADR2(\BU2/U0/N50778 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014_SW0 .INIT = 8'h75;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .O(\BU2/U0/N50778 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000820 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000820  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET ),
    .O(\BU2/U0/CHOICE2701 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>16 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/CHOICE1713 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455_128 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455_128  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0171 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR3(\BU2/U0/N51594 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2> .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/N51052 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>_SW0 .INIT = 8'h95;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [0]),
    .O(\BU2/U0/N51052 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .O(\BU2/U0/N51594 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193_129 .INIT = 16'h0203;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193_129  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR3(\BU2/U0/N50196 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193_SW0 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ),
    .O(\BU2/U0/N50196 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149_130 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149_130  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR3(\BU2/U0/N50568 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .O(\BU2/U0/N50568 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215571 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215571  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21559 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<3> .INIT = 16'hD0F2;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<3>  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .ADR2(\BU2/U0/N65648 ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<3>_SW1 .INIT = 16'hAAA9;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<3>_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [1]),
    .O(\BU2/U0/N65648 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<10>_rt_131 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<10>_rt_131  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [10]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<10>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>122 .INIT = 16'h8B00;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>122  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/CHOICE1790 ),
    .O(\BU2/U0/CHOICE1791 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n028723 .INIT = 16'h0888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n028723  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/N66126 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE ),
    .O(\BU2/U0/CHOICE2785 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0068_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX__n0068_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD ),
    .O(\BU2/U0/N53563 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt_132 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt_132  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21 .INIT = 8'h90;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>21  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .ADR2(\BU2/U0/CHOICE1713 ),
    .O(\BU2/U0/CHOICE1714 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt_133 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt_133  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt_134 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt_134  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_Mmux_BAD_FRAME_OUT_Result .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_Mmux_BAD_FRAME_OUT_Result  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ),
    .ADR2(\BU2/U0/N50165 ),
    .ADR3(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_COMB )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_Mmux_BAD_FRAME_OUT_Result_SW0 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_RX_Mmux_BAD_FRAME_OUT_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT ),
    .O(\BU2/U0/N50165 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt_135 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt_135  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0061_Result_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0061_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0297 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .O(\BU2/U0/N65965 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt_136 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt_136  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [9]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179_137 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179_137  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR3(\BU2/U0/N50537 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179_SW0 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .O(\BU2/U0/N50537 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<3> .INIT = 16'h0009;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<3>  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .ADR1(\BU2/U0/N65804 ),
    .ADR2(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR3(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<3>_SW1 .INIT = 8'h7F;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<3>_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .O(\BU2/U0/N65804 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125 .INIT = 16'h0027;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR1(\BU2/U0/N65986 ),
    .ADR2(\BU2/U0/N65984 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/CHOICE2752 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0060_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0060_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65784 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0060 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>109  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/CHOICE1738 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060_138 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060_138  (
    .ADR0(\BU2/U0/N65902 ),
    .ADR1(\BU2/U0/N65432 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .ADR3(\BU2/U0/CHOICE2587 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW12 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW12  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ),
    .ADR1(\BU2/U0/CHOICE1339 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .O(\BU2/U0/CHOICE1874 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010_139 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010_139  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .ADR3(\BU2/U0/N50134 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010_SW0 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT [0]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N50134 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mxor__n0014_Result1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mxor__n0014_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG_140 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG_140  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG_141 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG_141  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0007 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE_142 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE_142 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE_142  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4366 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt_143 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt_143  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<0>1 .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4370 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<0>1 .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n00071 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n00071  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0007 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04681 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04681  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4354 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<1>1 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>207 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>207  (
    .ADR0(\BU2/U0/CHOICE1820 ),
    .ADR1(\BU2/U0/CHOICE1831 ),
    .ADR2(\BU2/U0/CHOICE1845 ),
    .ADR3(\BU2/U0/CHOICE1863 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<5>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<1>1 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [1])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4366 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [4])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4362 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002<1>1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4366 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4354 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4358 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mxor__n0016_Result1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mxor__n0016_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0016 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4358 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4362 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<6>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002<1>1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000926 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000926  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME ),
    .ADR3(\BU2/U0/CHOICE2403 ),
    .O(\BU2/U0/CHOICE2404 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE_144 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE_144  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Ker229021 .INIT = 16'h000E;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Ker229021  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22904 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q [0]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C5 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C4 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C3 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C2 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TC ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C5 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C4 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C3 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C2 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TC ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C5 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C4 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C3 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C2 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TC ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C5 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C4 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C3 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C2 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TC ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF6  (
    .I(\BU2/U0/address_valid_early ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6q ),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5q ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TC_ASSIGN_I0 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI ),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_Q0_ASSIGN_LI_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_TQ0 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5q ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TC )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int3q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int2q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_FF1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1 ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int1q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [3]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ0 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_C1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TQ1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4362 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR_145 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR_145  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0009 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR_146 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR_146  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0008 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN_147 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN_147  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0007 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH_148 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH_148  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0024 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME_149 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME_149  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0005 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR_150 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR_150  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0018 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT_151 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT_151  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0013 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR_152 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR_152  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_2  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4293 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0022 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_153 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_153  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0019 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_N4870 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR_154 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR_154  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0011 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00051 .INIT = 16'h7770;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00051  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0005 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00071 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00071  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0007 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000965 .INIT = 16'hF800;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000965  (
    .ADR0(\BU2/U0/CHOICE2394 ),
    .ADR1(\BU2/U0/CHOICE2404 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR ),
    .ADR3(\BU2/U0/CHOICE2409 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0009 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060_SW1 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .O(\BU2/U0/N65902 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00111 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00111  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0023 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0011 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [5]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65516 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00131 .INIT = 16'h00AE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00131  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_ALIGNMENT_ERR_RD [0]),
    .ADR2(corehassgmii),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0013 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Ker165281 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Ker165281  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16530 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt_155 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt_155  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000894 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000894  (
    .ADR0(\BU2/U0/CHOICE2706 ),
    .ADR1(\BU2/U0/CHOICE2709 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0008 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Ker165331 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Ker165331  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16535 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00181 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00181  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0018 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00191 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n00191  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0019 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME_156 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME_156  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0015 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME_157 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME_157  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt_158 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt_158  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID_159 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID_159  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N16535 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022_Mxor__n0002_Result1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022_Mxor__n0002_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022__n0002 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_0  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4287 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR_160 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR_160  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0012 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut5 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut5  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4299 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_3  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4296 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo3 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut4 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut4  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4296 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut2 .INIT = 8'h18;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut2  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4290 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_1  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4290 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo2 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW12 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW12  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .ADR2(\BU2/U0/CHOICE1339 ),
    .O(\BU2/U0/CHOICE1866 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_norlut .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_norlut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4281 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut6 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut6  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4302 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_4  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4299 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_norcy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4281 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_nor_cyo )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_5  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4302 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo5 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut .INIT = 8'h81;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4284 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_ClkEn_INV1 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_ClkEn_INV1  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR_N4870 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut7 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut7  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4305 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_nor_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4284 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut1 .INIT = 8'h81;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [4]),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4287 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0059_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0059_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0296 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .O(\BU2/U0/N65780 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagecy_rn_6  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stage_cyo5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4305 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0023 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_34_161  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_34 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_37 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_34 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_38_162  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_37 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_34 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_38 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_331 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_331  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_33 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_33_163  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_33 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_36 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_33 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_37_164  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_36 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_33 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_37 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>7 .INIT = 16'h0604;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>7  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [0]),
    .O(\BU2/U0/CHOICE2716 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_32_165  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_32 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_35 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_32 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_36_166  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_35 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_32 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_36 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_311 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_311  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_31 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_31_167  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_31 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_34 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_31 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_35_168  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_34 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_31 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_35 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0114_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0114_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0114_Xo [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_30_169  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_30 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_33 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_30 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_34_170  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_33 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_30 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_34 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_291 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_291  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_29 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_29_171  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_29 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_32 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_29 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_33_172  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_32 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_29 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_33 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_32_173  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_32 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44_174 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44_174  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_43 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43_175 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43_175  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_42 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41_176 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41_176  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_40 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<9>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [9])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<9>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<9>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<9>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [8])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<8>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<7>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<7>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<6>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<6>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<5>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<5>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<4>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<4>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<3>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<3>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<2>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<1>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result43_G .INIT = 16'hB8BB;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RX_ER_Result43_G  (
    .ADR0(phyemacrxer),
    .ADR1(corehassgmii),
    .ADR2(\BU2/U0/CHOICE2628 ),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N66049 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>cy  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4255 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<0>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4255 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut29 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut29  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [10]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4252 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_27  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo21 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4249 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo22 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut28 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut28  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [9]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4249 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_26  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo20 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4246 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo21 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut27 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut27  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4246 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_25  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo19 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4243 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo20 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut26 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut26  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4243 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_24  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo18 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4240 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo19 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut25 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut25  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4240 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_23  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4237 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo18 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut24 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut24  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4237 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut23 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut23  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [22]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [23]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4234 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_21  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo16 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4231 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo17 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut22 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut22  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [20]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [21]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4231 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_20  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo15 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4228 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo16 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut21 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut21  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [18]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [19]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4228 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_19  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4225 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo15 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut20 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut20  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [16]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [17]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4225 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut19 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut19  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [31]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4222 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_17  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo13 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4219 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo14 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut18 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut18  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4219 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_16  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo12 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4216 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo13 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut17 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut17  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [27]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4216 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_15  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4213 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo12 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut16 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut16  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [25]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4213 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut15 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut15  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4210 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_13  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo10 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4207 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo11 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut14 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut14  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4207 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_12  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo9 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4204 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo10 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut13 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut13  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4204 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_11  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4201 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo9 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut12 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut12  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4201 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut11 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut11  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [38]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [39]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4198 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_9  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo7 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4195 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo8 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut10 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut10  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [36]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [37]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4195 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_8  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo6 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4192 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo7 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut9 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut9  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [34]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [35]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4192 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_7  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4189 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo6 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut8 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut8  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [32]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [33]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4189 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut7 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut7  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [15]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4186 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_5  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo4 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4183 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo5 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut6 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut6  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [12]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [13]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4183 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_4  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo3 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4180 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo4 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut5 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut5  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [10]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [11]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4180 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_3  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4177 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo3 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut4 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut4  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [9]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4177 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39_177 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39_177  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_38 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut3 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut3  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [46]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [47]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4172 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_1  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo1 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4169 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo2 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut2 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut2  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [44]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [45]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4169 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_0  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4166 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut1 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [42]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [43]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4166 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4163 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagelut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [40]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [41]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4163 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_35_178  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_35 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_38 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_35 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID_179 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID_179  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0052 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS_180 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS_180  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0051 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS_181 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS_181  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0050 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME_182 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME_182  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0104 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE_183 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE_183  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0047 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO_184 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO_184  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0046 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256_185 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256_185  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH_186 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH_186  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0110 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0161 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0042 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0041 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0040 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0039 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0038 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0037 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0036 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0035 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0034 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0033 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0032 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0149 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0024 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0023 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0022 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [2]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0030 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [3]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0029 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [4]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0028 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [5]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0027 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [6]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0026 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [7]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0024 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [8]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0023 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [9]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0022 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE [10]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE_187 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE_187  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_22  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo17 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4234 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0095 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_18  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo14 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4222 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0096 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET_188 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET_188  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0054 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0056 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0055 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0057 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0058 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0059 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0060 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0061 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0062 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0055 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0063 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0064 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0065 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0066 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0067 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH_189 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH_189  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE_190 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE_190  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0070 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0175 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT_191 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT_191  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00201 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00201  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0020 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00231 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00231  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0023 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00241 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00241  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0024 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00261 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00261  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0026 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00271 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00271  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0027 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00281 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00281  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0028 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00291 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00291  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0029 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00301 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00301  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0030 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00421 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00421  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0042 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00321 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00321  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0032 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00331 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00331  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0033 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00341 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00341  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0034 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00351 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00351  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0035 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00361 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00361  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0036 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00371 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00371  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0037 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00381 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00381  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0038 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00391 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00391  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0039 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00401 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00401  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0040 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00411 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00411  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0041 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0045_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0045_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [12]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0045 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161201 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker161201  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_192 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_192  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00501 .INIT = 16'h7770;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00501  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0050 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>62 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<5>62  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [13]),
    .O(\BU2/U0/CHOICE3038 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n001236 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n001236  (
    .ADR0(\BU2/U0/CHOICE2595 ),
    .ADR1(\BU2/U0/CHOICE2600 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00551 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00551  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0055 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In_193 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In_193  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER ),
    .ADR2(\BU2/U0/N57873 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00621 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00621  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0098 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0062 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00631 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00631  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0097 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0063 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00641 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00641  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0096 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0064 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00651 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00651  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0095 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0065 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00661 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00661  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0094 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0066 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00671 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00671  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0093 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0067 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00441 .INIT = 16'h2276;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n00441  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0044 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_G .INIT = 16'h1D3C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>80_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/N66054 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00731 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00731  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00751 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00751  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0075 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448_194 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448_194  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR3(\BU2/U0/N50513 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0116_Xo<0>1 .INIT = 8'h69;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0116_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0116_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0165 ),
    .O(\BU2/U0/N50513 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_42_195  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_42 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_45 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_42 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_46_196  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_45 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_42 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_46 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_43_197  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_42 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_39 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_43 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_11 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_11  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker160901 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker160901  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16092 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_39_198  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_39 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_42 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_39 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_40_199  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_40 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_43 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_40 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42_200 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42_200  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_41 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In_SW0 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .O(\BU2/U0/N57873 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38_201 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38_201  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_37 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01761 .INIT = 8'h8F;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01761  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01101 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01101  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0103 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0110 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_41_202  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_40 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_37 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_41 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_351 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_351  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_35 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40_203 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40_203  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_39 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_40_204  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_39 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_36 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_40 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_43_205  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_43 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_46 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_43 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_36_206  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_36 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_39 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_36 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30_207 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30_207  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_29 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31_208 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31_208  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_30 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_01 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_01  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_0 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_37_209  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_37 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_40 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_37 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_41 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_41  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_41_210  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_41 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_44 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_41 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_42_211  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_41 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_38 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_42 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32_212 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32_212  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_31 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_38_213  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_38 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_41 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_38 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33_214 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33_214  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_32 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_51 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_51  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_5 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_21 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_21  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_2 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34_215 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34_215  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_33 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01881 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01881  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35_216 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35_216  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_34 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36_217 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36_217  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_35 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_44_218  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_43 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_40 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_44 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37_219 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37_219  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_sum_36 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0176 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_31 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_31  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_3 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0059_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0059_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65780 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0059 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt_220 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt_220  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01611 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01611  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0161 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW18 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014_SW18  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/CHOICE1878 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01751 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01751  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0175 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01811 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01811  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0181 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0073 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG_221 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG_221  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH_222 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH_222  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0075 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0179 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME_223 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME_223  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME_224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME_224  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0077 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0181 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0078 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0079 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0080 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0081 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0082 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH_225 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH_225  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME_226 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME_226  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0084 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16122 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT_227 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT_227  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0086 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0188 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_228 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_228  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker160851 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Ker160851  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16087 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05121 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05121  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0512 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_361 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_361  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_36 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Mmux__n0052_Result1 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Mmux__n0052_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16087 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0052 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<10>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<10>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DECODE_FRAME__n0000<9>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0000 [10])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_14  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo11 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4210 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0093 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_10  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo8 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4198 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0097 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_6  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo5 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4186 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0094 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_2  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo2 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4172 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0098 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stagecy_rn_28  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_Eq_stage_cyo22 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N4252 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0103 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_45_229  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_44 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_41 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_45 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_39_230  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_38 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_35 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_cy_39 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME_231 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME_231  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0029 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00221 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00221  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0022 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00231 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00231  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0023 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00181 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00181  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0018 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00211 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00211  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0021 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00301 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00301  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0030 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE_232 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE_232  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0030 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0059 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>120 .INIT = 16'h9200;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>120  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .ADR3(\BU2/U0/CHOICE1738 ),
    .O(\BU2/U0/CHOICE1739 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00271 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00271  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0027 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00151 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00151  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0015 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0324_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [1]),
    .O(\BU2/U0/N53310 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD_233 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD_233  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0017 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA_234 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA_234  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0027 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00241 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00241  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0024 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0061_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0061_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N54124 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0061 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD_235 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD_235  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0014 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt_236 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt_236  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n00441 .INIT = 16'h2276;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n00441  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WREN_REG ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0044 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt_237 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt_237  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD_238 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD_238  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0015 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD_239 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD_239  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0018 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD_240 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD_240  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0060 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0021 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0022 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0023 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0024 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026 ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<1>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [33]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [41]),
    .O(\BU2/U0/CHOICE3067 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_3 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0062 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [3]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_4 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0061 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [4]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_5 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0060 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [5]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_31 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_31  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0034 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_30 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_30  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0035 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_29 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_29  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0036 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_28 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_28  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0037 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_7 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0058 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [7]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0131_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0131_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0317 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0132_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0132_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0133_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0133_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0318 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0134_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0134_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0135_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0135_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0136_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0136_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278<1>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0157_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0157_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0143_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0143_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0144_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0144_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0055_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0055_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0055 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_1 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0064 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [1]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0159_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0159_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0164_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0164_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0296 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0046_Result1 .INIT = 8'h6A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0046_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0046 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0166_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0166_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0297 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0170_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0170_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0299 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>59 .INIT = 16'h1800;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<1>59  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .ADR3(\BU2/U0/CHOICE1830 ),
    .O(\BU2/U0/CHOICE1831 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_10 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_10  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0055 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [10]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_13 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_13  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0052 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [13]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_12 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_12  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0053 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [12]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_15 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_15  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0050 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [15]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_14 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_14  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0051 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [14]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_17 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_17  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0048 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [17]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_16 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_16  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0049 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [16]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_19 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_19  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0046 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [19]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_18 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_18  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0047 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [18]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_9 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_9  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0056 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [9]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_6 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0059 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [6]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_21 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_21  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0044 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [21]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_20 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_20  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0045 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [20]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_23 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_23  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0042 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [23]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_22 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_22  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0043 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [22]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_25 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_25  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0040 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_24 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_24  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0041 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_27 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_27  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0038 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_26 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_26  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0039 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<13>161_G .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<13>161_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [7]),
    .O(\BU2/U0/N66059 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_0 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0065 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [0]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083_241 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083_241  (
    .ADR0(\BU2/U0/N65628 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_8 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0057 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [8]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0057_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0057_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0126_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0057 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0056_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0056_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0056 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<14>161_G .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<14>161_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [8]),
    .O(\BU2/U0/N66064 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_11 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_11  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0054 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [11]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0042_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0042_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [15]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0042 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0041_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0041_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [16]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0277 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0041 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0040_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0040_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [17]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0040 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0035_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0035_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [22]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0318 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0035 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083_SW1 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0083_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD ),
    .O(\BU2/U0/N65628 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0034_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0034_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [23]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0034 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0043_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0043_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0043 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0054_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0054_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [24]),
    .O(\BU2/U0/N65938 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0054_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0054_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [3]),
    .ADR1(\BU2/U0/N65938 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0295 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0054 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0061_Result_SW0 .INIT = 8'h69;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0061_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0297 [2]),
    .O(\BU2/U0/N54124 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0051_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0051_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0116_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0051 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0050_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0050_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/N65934 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0050_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0050_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [7]),
    .ADR1(\BU2/U0/N65934 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0050 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0113_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0113_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0113_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0049_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0049_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0114_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0049 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0112_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0112_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0112_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0048_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0048_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0113_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0048 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0101_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0101_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0101_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0047_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0047_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0112_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0047 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0039_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0039_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .O(\BU2/U0/N65930 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0039_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0039_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [18]),
    .ADR1(\BU2/U0/N65930 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0039 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0038_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0038_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [28]),
    .O(\BU2/U0/N65926 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0038_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0038_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [19]),
    .ADR1(\BU2/U0/N65926 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0277 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0038 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0037_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0037_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [20]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0317 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0037 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0114_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0114_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0114_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0036_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0036_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [21]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0319 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0101_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0036 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0118_Xo<3>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0118_Xo<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0316 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0294 [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0118_Xo [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0044_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0044_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [13]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0044 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0053_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0053_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0318 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0118_Xo [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0053 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0065_Result1 .INIT = 8'h72;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0065_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0278 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0065 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0137_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0137_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0277 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0052_Result1_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0052_Result1_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0117_Xo [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0102_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [29]),
    .O(\BU2/U0/N65776 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0052_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mmux__n0052_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [5]),
    .ADR1(\BU2/U0/N65776 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0320 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0052 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0045_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0045_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [12]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0045 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_24_242  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_24 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_26 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_24 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_27_243  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_26 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_24 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_27 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00441 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00441  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .ADR2(\BU2/U0/CHOICE1339 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_23_244  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_23 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_25 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_23 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_26_245  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_25 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_23 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_26 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_22_246  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_22 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_24 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_22 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_25_247  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_24 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_22 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_25 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_24_248  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/N66102 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_24 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_25_249  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_25 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_27 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_25 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG_250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG_250  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RX_DV ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_281 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_281  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_28 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_30_251  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_29 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_27 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_30 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC_252 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC_252  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n0006 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt_253 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt_253  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_29_254  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_28 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_26 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_29 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN<5>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN<5>1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(corehassgmii),
    .ADR2(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[5] )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00071 .INIT = 16'hFF7F;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00071  (
    .ADR0(\BU2/U0/CHOICE2494 ),
    .ADR1(\BU2/U0/CHOICE2501 ),
    .ADR2(\BU2/U0/CHOICE2486 ),
    .ADR3(\BU2/U0/N65358 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0007 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_26 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_26 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_26  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_26 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [4])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_25 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_25 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_25  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_25 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [3])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_23 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_23  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_23 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [1])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_22 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_22  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_22 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN<3>1 .INIT = 8'hBF;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN<3>1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(corehassgmii),
    .ADR2(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DIN[3] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_26_255  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_26 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_28 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_26 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_28_256  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_28 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_30 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_28 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_28 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_28 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_28  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_28 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [6])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_27 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_27 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_27  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_27 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [5])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_24 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_24 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_24  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_24 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [2])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_27_257  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_27 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_29 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_sum_27 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42  (
    .I(tieemacconfigvec_7[42]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [42]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41  (
    .I(tieemacconfigvec_7[41]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [41]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40  (
    .I(tieemacconfigvec_7[40]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [40]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39  (
    .I(tieemacconfigvec_7[39]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [39]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38  (
    .I(tieemacconfigvec_7[38]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [38]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37  (
    .I(tieemacconfigvec_7[37]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [37]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36  (
    .I(tieemacconfigvec_7[36]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [36]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35  (
    .I(tieemacconfigvec_7[35]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [35]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34  (
    .I(tieemacconfigvec_7[34]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [34]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33  (
    .I(tieemacconfigvec_7[33]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [33]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32  (
    .I(tieemacconfigvec_7[32]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [32]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31  (
    .I(tieemacconfigvec_7[31]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [31]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30  (
    .I(tieemacconfigvec_7[30]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [30]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29  (
    .I(tieemacconfigvec_7[29]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [29]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28  (
    .I(tieemacconfigvec_7[28]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [28]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27  (
    .I(tieemacconfigvec_7[27]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [27]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26  (
    .I(tieemacconfigvec_7[26]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [26]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25  (
    .I(tieemacconfigvec_7[25]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [25]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24  (
    .I(tieemacconfigvec_7[24]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [24]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23  (
    .I(tieemacconfigvec_7[23]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [23]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22  (
    .I(tieemacconfigvec_7[22]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [22]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21  (
    .I(tieemacconfigvec_7[21]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [21]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20  (
    .I(tieemacconfigvec_7[20]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [20]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19  (
    .I(tieemacconfigvec_7[19]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [19]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18  (
    .I(tieemacconfigvec_7[18]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [18]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17  (
    .I(tieemacconfigvec_7[17]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [17]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16  (
    .I(tieemacconfigvec_7[16]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [16]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15  (
    .I(tieemacconfigvec_7[15]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14  (
    .I(tieemacconfigvec_7[14]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13  (
    .I(tieemacconfigvec_7[13]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12  (
    .I(tieemacconfigvec_7[12]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11  (
    .I(tieemacconfigvec_7[11]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10  (
    .I(tieemacconfigvec_7[10]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9  (
    .I(tieemacconfigvec_7[9]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8  (
    .I(tieemacconfigvec_7[8]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7  (
    .I(tieemacconfigvec_7[7]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6  (
    .I(tieemacconfigvec_7[6]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5  (
    .I(tieemacconfigvec_7[5]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4  (
    .I(tieemacconfigvec_7[4]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3  (
    .I(tieemacconfigvec_7[3]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2  (
    .I(tieemacconfigvec_7[2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1  (
    .I(tieemacconfigvec_7[1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0  (
    .I(tieemacconfigvec_7[0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n00001 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n00011 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD_258 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD_258  (
    .I(tieemacconfigvec_7[63]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD_259 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD_259  (
    .I(tieemacconfigvec_7[48]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD_260 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD_260  (
    .I(tieemacconfigvec_7[51]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD_261 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD_261  (
    .I(tieemacconfigvec_7[49]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD_262 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD_262  (
    .I(tieemacconfigvec_7[52]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47  (
    .I(tieemacconfigvec_7[47]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [47]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG_263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG_263  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0030 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(NlwRenamedSig_OI_emacclientrxstats[0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(NlwRenamedSig_OI_emacclientrxstats[1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0029 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [3]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [4]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [5]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[10]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [6]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[11]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[12]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [8]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[13]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [9]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[14]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [10]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[15]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [11]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[16]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [12]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[17]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH [13]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[18]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[19]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[20]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[21]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[22]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_LENGTH_TYPE_ERROR ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[25]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0028 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstats_6[26]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG_264 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG_264  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Ker227431 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Ker227431  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22745 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxstatsvld),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CRC1000_EN_265 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_CRC1000_EN_265  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV100_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CRC1000_EN ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV100_REG_266 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV100_REG_266  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV100_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT_267 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT_267  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT_268 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT_268  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0025 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT_269 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT_269  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0024 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT_270 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT_270  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0023 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT_271 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT_271  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0022 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN_272 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN_272  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV10_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV10_REG_273 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV10_REG_273  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CLK_DIV10_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT_274 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT_274  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT_275 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT_275  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0019 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT_276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT_276  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0018 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT_277 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT_277  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0017 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT_278 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT_278  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0016 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR_279 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR_279  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_2 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0063 ),
    .SRST(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [2]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_341 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_341  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_34 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD_280 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD_280  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0016 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG_281 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG_281  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .SET(GND),
    .RST(GSR)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_28_282  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_27 ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_25 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_cy_28 )
  );
  X_AND2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int4q ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_TC ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int5 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8 [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_8  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [7]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [8]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG_283 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG_283  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0033 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG_284 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG_284  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0034 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WR_REG_285 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WR_REG_285  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WR_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD_286 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD_286  (
    .I(NlwRenamedSig_OI_speedis10100),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0001 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CRC_CE1 .INIT = 16'hB8BB;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_CRC_CE1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CRC1000_EN ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_CRC100_EN ),
    .ADR3(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CRC_CE )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4374 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43  (
    .I(tieemacconfigvec_7[43]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [43]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR_287 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR_287  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RX_DV ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WR_REG_288 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WR_REG_288  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WR_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR_289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR_289  (
    .I(\BU2/U0/TRIMAC_INST_INT_GMII_RX_ER ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1_290 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1_290  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RX_DV ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2_291 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2_291  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00161 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN__n00161  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0016 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00171 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00171  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0017 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44  (
    .I(tieemacconfigvec_7[44]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [44]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00191 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00191  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0019 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46  (
    .I(tieemacconfigvec_7[46]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [46]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>62 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>62  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [10]),
    .O(\BU2/U0/CHOICE3015 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00221 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN__n00221  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0022 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00231 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00231  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0023 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45  (
    .I(tieemacconfigvec_7[45]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RESET_CRC ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD [45]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00251 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00251  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0025 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4378 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001284 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001284  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .O(\BU2/U0/CHOICE2928 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00281 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN__n00281  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0028 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00291 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN__n00291  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0029 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00301 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN__n00301  (
    .ADR0(tieemacconfigvec_7[50]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_int6q ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0030 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6_292 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6_292  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG5 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>39_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>39_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [4]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(\BU2/U0/N65512 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00204 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00204  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [5]),
    .O(\BU2/U0/CHOICE2122 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7_293 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7_293  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<2>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [10]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<3>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[3]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [11]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<1>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<1>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [9]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<0>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<0>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [8]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00181 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00181  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0018 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n00241 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN__n00241  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0024 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW15 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015_SW15  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_FORCE_QUIET ),
    .O(\BU2/U0/CHOICE1868 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .WRITE_MODE_A = "READ_FIRST";
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_A = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .INIT_B = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .SRVAL_A = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0 .SRVAL_B = 36'h000000000;
  X_RAMB16_S36_S36 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0  (
    .CLKA(rxgmiimiiclk),
    .CLKB(rxcoreclk),
    .ENA(\BU2/U0/address_valid_early ),
    .ENB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .SSRA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SSRB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .WEA(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .WEB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .GSR(GSR),
    .ADDRA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]}),
    .ADDRB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]}),
    .DIA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_ER_WR_REG , \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WR_REG , \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [8], 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [7], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [6], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [5], 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [4], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [3], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [2], 
\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [1], \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [0]}),
    .DIB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DIPA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DIPB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DOA({\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[31]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[30]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[29]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[28]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[27]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[26]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[25]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[24]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[23]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[22]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[21]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[20]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[19]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[18]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[17]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[16]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[15]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[14]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[13]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[12]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[11]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[10]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[9]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[8]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[7]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[6]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[5]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[4]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOA[0]_UNCONNECTED }),
    .DOPA({\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPA[0]_UNCONNECTED }),
    .DOB({\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[31]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[30]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[29]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[28]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[27]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[26]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[25]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[24]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[23]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[22]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[21]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[20]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[19]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[18]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[17]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[16]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[15]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[14]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[13]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[12]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOB[11]_UNCONNECTED , \BU2/U0/TRIMAC_INST_RXGEN__n0108 [1], 
\BU2/U0/TRIMAC_INST_RXGEN__n0106 [1], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [15], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [14], 
\BU2/U0/TRIMAC_INST_RXGEN__n0109 [13], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [12], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [11], 
\BU2/U0/TRIMAC_INST_RXGEN__n0109 [10], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [9], \BU2/U0/TRIMAC_INST_RXGEN__n0109 [8], 
\BU2/U0/TRIMAC_INST_RXGEN_RXD_ALIGNMENT_ERR_RD [0]}),
    .DOPB({\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mram_mem_inst_ramb_0_DOPB[0]_UNCONNECTED })
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<5>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<5>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [13]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [5])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<7>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[7]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [15]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [7])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1_294 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1_294  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RX_ERR ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6_295 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6_295  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG5 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7_296 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7_296  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<4>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<4>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[4]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [12]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [4])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [7]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00061 .INIT = 16'h00F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00061  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxdv),
    .ADR2(\BU2/U0/CHOICE1120 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n0006 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<6>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RXD_Result<6>1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0109 [14]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RXD [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04545 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04545  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .O(\BU2/U0/CHOICE2651 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID_297 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID_297  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RX_ERR_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RX_ERR_Result1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxer),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0108 [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RX_ERR )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [2]),
    .RST(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4370 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4378 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [0]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [0]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [1]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [1]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [2]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [2]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [3]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4370 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046181 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046181  (
    .ADR0(\BU2/U0/CHOICE3153 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/CHOICE3145 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0461 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [3]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [4]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [4]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [5]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [5]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [6]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [6]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [7]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0000 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4354 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4366 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [4])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [0])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4362 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012186 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012186  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [1]),
    .ADR2(\BU2/U0/CHOICE3193 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022_Mxor__n0002_Result1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022_Mxor__n0002_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Msub__n0022__n0002 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker227431 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Ker227431  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22745 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG_298 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG_298  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WREN_REG ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [7]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [8]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WR_REG_299 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WR_REG_299  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WR_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WR_REG_300 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WR_REG_300  (
    .I(\BU2/U0/N66295 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WR_REG ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .WRITE_MODE_A = "READ_FIRST";
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_A = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .INIT_B = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .SRVAL_A = 36'h000000000;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0 .SRVAL_B = 36'h000000000;
  X_RAMB16_S36_S36 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0  (
    .CLKA(txcoreclk),
    .CLKB(txgmiimiiclk),
    .ENA(\BU2/U0/address_valid_early ),
    .ENB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .SSRA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SSRB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .WEA(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .WEB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .GSR(GSR),
    .ADDRA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]}),
    .ADDRB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]}),
    .DIA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WR_REG , \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_EN_WR_REG , \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [8], 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [7], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [6], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [5], 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [4], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [3], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [2], 
\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [1], \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_D_WR_REG [0]}),
    .DIB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DIPA({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DIPB({\NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , \NlwRenamedSig_OI_BU2/emacphymclkout , 
\NlwRenamedSig_OI_BU2/emacphymclkout }),
    .DOA({\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[31]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[30]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[29]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[28]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[27]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[26]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[25]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[24]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[23]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[22]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[21]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[20]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[19]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[18]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[17]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[16]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[15]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[14]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[13]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[12]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[11]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[10]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[9]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[8]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[7]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[6]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[5]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[4]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOA[0]_UNCONNECTED }),
    .DOPA({\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPA[0]_UNCONNECTED }),
    .DOB({\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[31]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[30]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[29]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[28]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[27]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[26]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[25]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[24]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[23]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[22]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[21]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[20]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[19]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[18]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[17]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[16]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[15]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[14]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[13]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[12]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOB[11]_UNCONNECTED , \BU2/U0/TRIMAC_INST_TXGEN__n0038 [1], 
\BU2/U0/TRIMAC_INST_TXGEN__n0037 [1], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [15], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [14], 
\BU2/U0/TRIMAC_INST_TXGEN__n0035 [13], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [12], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [11], 
\BU2/U0/TRIMAC_INST_TXGEN__n0035 [10], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [9], \BU2/U0/TRIMAC_INST_TXGEN__n0035 [8], 
\BU2/U0/TRIMAC_INST_TXGEN__n0039 [1]}),
    .DOPB({\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[3]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[2]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[1]_UNCONNECTED , 
\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mram_mem_inst_ramb_0_DOPB[0]_UNCONNECTED })
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt_301 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt_301  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC4_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0014 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0016 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [0]),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4358 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [2])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4354 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [1])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4378 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [7])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4374 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4374 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0116_Xo<0>1 .INIT = 8'h69;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0116_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0116_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<12>161_G .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<12>161_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [6]),
    .O(\BU2/U0/N66069 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2> .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/N50978 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [2])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mxor__n0014_Result1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mxor__n0014_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG_302 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG_302  (
    .I(\BU2/U0/N66129 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_ER_WREN_REG ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG_303 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG_303  (
    .I(\BU2/U0/N66231 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0001 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE_304 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE_304 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE_304  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0010 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4366 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<0>1 .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4370 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<0>1 .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RX_DV_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_Mmux_INT_RX_DV_Result1  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxdv),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0106 [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_INT_RX_DV )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4354 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<1>1 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>207 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>207  (
    .ADR0(\BU2/U0/CHOICE1714 ),
    .ADR1(\BU2/U0/CHOICE1725 ),
    .ADR2(\BU2/U0/CHOICE1739 ),
    .ADR3(\BU2/U0/CHOICE1757 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_OCCUPANCY [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<1>1 .INIT = 16'hA8AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0000 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4362 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR__n0004 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002<1>1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR__n0002 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4366 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0__n00001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4358 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mxor__n0016_Result1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mxor__n0016_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0016 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4358 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4362 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002<1>1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR__n0002 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n004531 .INIT = 16'hE0FF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n004531  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_N22904 ),
    .ADR2(\BU2/U0/CHOICE3250 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0007 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0045 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE_305 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE_305  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n0012 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5_306 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5_306  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5-In ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt_307 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt_307  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>_SW0 .INIT = 8'h95;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [0]),
    .O(\BU2/U0/N50978 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5-In1 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5-In1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_N21825 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5-In )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [2]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<0>1 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<1>1 .INIT = 8'h09;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<2>1 .INIT = 16'hEEEB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1_308 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1_308  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [3]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [3]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2_309 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2_309  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4354 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT__n0001 [0]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT [0]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt_310 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt_310  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004510 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004510  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [7]),
    .O(\BU2/U0/CHOICE2540 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791_SW0 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01791_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .O(\BU2/U0/N65254 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3_311 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3_311  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_Ker218231 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_Ker218231  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS ),
    .ADR1(tieemacconfigvec_7[55]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_N21825 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_31 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_31  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0034 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_30 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_30  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0035 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_29 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_29  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0036 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_28 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_28  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0037 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_7 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0058 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [7]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0131_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0131_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0317 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0132_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0132_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0133_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0133_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0318 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0134_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0134_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0135_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0135_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0136_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0136_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278<1>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0159_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0159_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0143_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0143_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0144_Result1 .INIT = 4'h9;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0144_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0055_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0055_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0294 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0055 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_1 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0064 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [1]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_FORCE_QUIET_Result16_G .INIT = 16'h000E;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_FORCE_QUIET_Result16_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .O(\BU2/U0/N66074 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0164_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0164_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0296 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0046_Result1 .INIT = 8'h6A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0046_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0046 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0166_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0166_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0297 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0170_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0170_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0299 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN_312 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN_312  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21490 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [0]),
    .ADR3(\BU2/U0/N53396 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_10 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0055 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [10]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_13 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0052 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [13]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_12 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0053 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [12]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_15 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_15  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0050 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [15]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_14 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0051 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [14]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_17 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_17  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0048 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [17]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_16 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_16  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0049 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [16]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_19 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_19  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0046 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [19]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_18 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_18  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0047 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [18]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_9 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0056 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [9]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_6 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0059 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [6]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_21 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_21  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0044 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [21]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_20 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_20  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0045 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [20]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_23 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_23  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0042 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [23]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_22 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_22  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0043 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [22]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_25 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_25  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0040 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_24 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_24  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0041 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_27 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_27  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0038 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_26 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_26  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0039 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_301 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_301  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_30 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_0 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0065 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [0]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>162 .INIT = 16'h01D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<2>162  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [2]),
    .O(\BU2/U0/CHOICE1698 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_8 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0057 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [8]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0057_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0057_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0126_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0057 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0056_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0056_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0294 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0056 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036_313 .INIT = 16'h5455;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036_313  (
    .ADR0(\BU2/U0/N65906 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .ADR2(\BU2/U0/N65432 ),
    .ADR3(\BU2/U0/CHOICE2587 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_11 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0054 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [11]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0042_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0042_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [15]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0042 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0041_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0041_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [16]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0277 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0041 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0040_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0040_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [17]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0040 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0035_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0035_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [22]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0318 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0035 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0157_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0157_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0294 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036_SW1 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0036_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .O(\BU2/U0/N65906 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0034_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0034_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [23]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0034 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0045 .INIT = 16'h222A;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0045  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [3]),
    .ADR1(\BU2/U0/N52548 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0043_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0043_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0043 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0054_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0054_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/N65922 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0054_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0054_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [3]),
    .ADR1(\BU2/U0/N65922 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0054 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>161_G .INIT = 16'hAAFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>161_G  (
    .ADR0(\BU2/U0/CHOICE1945 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .O(\BU2/U0/N66079 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0051_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0051_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0116_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0051 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0050_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0050_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/N65918 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0050_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0050_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [7]),
    .ADR1(\BU2/U0/N65918 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0050 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0113_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0113_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0113_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0049_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0049_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0114_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0049 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0112_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0112_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0112_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0048_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0048_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [9]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0113_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0048 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0101_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0101_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0101_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0047_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0047_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0112_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0047 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0039_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0039_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/N65914 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0039_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0039_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [18]),
    .ADR1(\BU2/U0/N65914 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0039 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0038_Result1_SW1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0038_Result1_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .O(\BU2/U0/N65910 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0038_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0038_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [19]),
    .ADR1(\BU2/U0/N65910 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0277 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0038 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo<0>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0037_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0037_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [20]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0317 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0037 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0137_Result1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_Mxor__n0137_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [25]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK_REG [31]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FCS_CHECK__n0277 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0036_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0036_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [21]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0101_Xo [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0036 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0118_Xo<3>1 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0118_Xo<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0294 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0118_Xo [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0044_Result1 .INIT = 16'h6CC6;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0044_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [13]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0044 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0053_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0053_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0318 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0118_Xo [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0053 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0065_Result1 .INIT = 8'h72;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0065_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0278 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0065 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0058_Result_SW0 .INIT = 16'h6996;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0058_Result_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0317 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0316 [1]),
    .O(\BU2/U0/N53888 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0052_Result1_SW0 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0052_Result1_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0117_Xo [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mxor__n0102_Xo [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .O(\BU2/U0/N65772 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0052_Result1 .INIT = 16'h96AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0052_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [5]),
    .ADR1(\BU2/U0/N65772 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0052 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0038_Result1 .INIT = 16'h1F0E;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0038_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .ADR2(tieemacconfigvec_7[66]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0038 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4335 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4335 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4335 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4331 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4331 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4331 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4327 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4327 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4327 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4323 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4323 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4323 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4319 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4319 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4319 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4315 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4315 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4315 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [0])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0045_SW0 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n0045_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/N52548 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [6]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4343 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088 [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [15]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [14]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [13]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [12]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [11]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [10]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [9]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [8]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [8]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [7]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [6]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [5]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [4]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [3]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [2]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [17]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [17]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [18]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [18]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[4]),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [1]),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[5] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0_314 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0_314  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1_315 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1_315  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2_316 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2_316  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3_317 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3_317  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt_318 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt_318  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n001213 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n001213  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .ADR2(\BU2/U0/CHOICE2590 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .O(\BU2/U0/CHOICE2595 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0100 [3]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX [2]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4_319 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4_319  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[6] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[7] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[8] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4339 ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4339 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [11]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4339 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<8>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_LPM_COUNTER_7__n0002<8>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_N4343 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [8]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [2]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker212881 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker212881  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21290 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026_320 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026_320  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .ADR3(\BU2/U0/N50462 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n00001 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .ADR2(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [0]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [0]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026_SW0 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0026_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ),
    .O(\BU2/U0/N50462 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03861 .INIT = 16'hBBB0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03861  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001284 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001284  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [2]),
    .O(\BU2/U0/CHOICE3181 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN_SW0 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [11]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [3]),
    .O(\BU2/U0/N53396 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0058_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0058_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0319 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N53888 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0058 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03131 .INIT = 16'h3B08;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03131  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21290 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0313 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01561 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01561  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_ACK_IN )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215231 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker215231  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<2>1 .INIT = 16'hABA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [12]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_11__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [11]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [10]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_9__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [9]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_8__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [8]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_7__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [7]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_6__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [6]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_5__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [5]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [4]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21559 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [3]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_2__n0000 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [2]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [1]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [0]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [13]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21559 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [14]),
    .CE(VCC)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001023_SW0 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001023_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR ),
    .O(\BU2/U0/N65436 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000824 .INIT = 16'hFF8A;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000824  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH ),
    .ADR3(\BU2/U0/CHOICE2701 ),
    .O(\BU2/U0/CHOICE2702 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [6]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_64_321  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_64 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_69 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_64 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10_322 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10_322  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [8]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5_323 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5_323  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[9] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[10] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[10]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[11] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[11]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51_324 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51_324  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_50 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[12] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[12]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[13] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[13]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<6>1 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [25]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52_325 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52_325  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_51 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[14] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[14]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[15] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[15]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n00011 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .ADR2(tieemacconfigvec_7[66]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0001 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW__n00091 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW__n00091  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ),
    .ADR3(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(emacclientrxstats_6[23])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut71 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut71  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4625 ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_5  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo5 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4622 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo6 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut6 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut6  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64 ),
    .ADR3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4622 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_4  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo4 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4619 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo5 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut5 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut5  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62 ),
    .ADR3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4619 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_3  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo3 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4616 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo4 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut4 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut4  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .ADR3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4616 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_2  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo2 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4613 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo3 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut3 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut3  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58 ),
    .ADR3(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4613 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_1  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4610 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo2 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut2 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut2  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56 ),
    .ADR3(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4610 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_0  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4607 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo1 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut1 .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4607 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4604 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut .INIT = 16'h9009;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagelut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52 ),
    .ADR3(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4604 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[16] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[16]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4600 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4596 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4596 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4596 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4592 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4592 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4592 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4588 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4588 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4588 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<11>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<3>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0537<10>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2_326 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2_326  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<16>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[17] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[15] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[14] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<14>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[13] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<13>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[12] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<12>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[11] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<2>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<11>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4566 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[10] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4566 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<10>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046173 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046173  (
    .ADR0(\BU2/U0/N65408 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/CHOICE3153 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>cy  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4562 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<9>_cyo )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[8] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[6] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<6>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[5] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<5>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<5>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[4] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<4>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<4>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[3] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<3>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<3>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4548 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[2] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4548 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<2>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[1] )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_IFG_DELAY_HELD<1>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001248 .INIT = 16'h9D80;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001248  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .O(\BU2/U0/CHOICE2918 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>cy  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4542 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[17] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[17]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<18>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<18>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [18]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4538 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4534 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [17])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4534 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [17]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4534 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4530 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [16])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4530 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<16>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [16]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4530 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4526 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [15])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4526 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<15>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [15]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4526 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4522 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [14])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4522 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<14>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [14]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4522 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4518 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [13])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4518 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<13>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4514 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [12])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4514 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<12>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4510 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [11])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4510 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<11>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4506 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [10])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4506 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<10>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4502 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [9])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4502 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<9>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4498 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [8])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4498 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<8>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4494 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4494 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<7>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4490 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4490 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<6>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4486 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4486 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<5>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4482 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4482 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<4>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4478 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4478 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<3>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4474 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4474 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<2>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4470 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4470 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<1>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [0])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[18] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[18]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [8])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<8>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<8>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<7>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<7>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<6>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<5>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<4>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<3>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<2>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<2>_cyo )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<1>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt_327 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt_327  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q7_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>cy  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4446 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<0>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4446 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[19]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<14>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<14>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [14]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4442 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4438 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [13])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4438 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [13]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4438 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4434 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [12])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4434 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<12>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [12]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4434 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4430 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [11])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4430 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<11>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [11]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4430 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4426 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [10])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4426 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<10>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [10]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4426 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4422 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [9])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4422 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<9>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4422 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4418 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [8])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4418 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<8>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4418 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4414 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4414 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4414 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4410 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4410 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4410 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4406 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4406 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4406 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4402 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4402 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4402 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4398 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4398 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4398 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4394 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4394 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4394 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4390 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4390 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4390 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [0])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_STATUS_VALID ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID.GSR.OR ),
    .CLK(txcoreclk),
    .O(NlwRenamedSig_OI_emacclienttxstatsvld),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[20]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE_328 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE_328  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0530 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED_329 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED_329  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0146 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0528 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2_330 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2_330  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0144 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0527 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2 ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET_331 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET_331  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0202 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0526 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS_332 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS_332  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID_333 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID_333  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION_334 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION_334  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0525 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS_335 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS_335  (
    .I(\BU2/U0/N66290 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0524 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [3]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [3]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT_336 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT_336  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0523 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH_337 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH_337  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[21]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[22]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14_338 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14_338  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN_339 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN_339  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_VLAN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL_340 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL_340  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_CONTROL ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH_341 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH_341  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0132 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH_342 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH_342  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH_343 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH_343  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0132 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH_344 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH_344  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0131 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH_345 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH_345  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0130 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH_346 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH_346  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0129 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH_347 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH_347  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0128 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS_348 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS_348  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0200 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0514 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2_349 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2_349  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0123 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0513 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN_350 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN_350  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0123 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0512 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID_351 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID_351  (
    .I(\BU2/U0/N66193 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0511 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL_352 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL_352  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0198 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT_353 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT_353  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0197 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START_354 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START_354  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0196 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0510 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX_355 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX_355  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0115 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [8]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [9]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [10]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [10]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [11]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [11]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [12]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [12]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7_356 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7_356  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7_357 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7_357  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7_358 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7_358  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7_359 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7_359  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7_360 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7_360  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE_361 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE_361  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0111 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION_362 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION_362  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0193 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_363 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_363  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0192 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_364 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_364  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0191 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_365 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_365  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0190 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_366 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_366  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_367 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_367  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0189 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_368 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_368  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0188 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY_369 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY_369  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0104 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0475 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN_370 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN_370  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0474 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[23]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED_371 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED_371  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0186 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0473 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED_372 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED_372  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0472 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED_373 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED_373  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0095 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0471 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63_374 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63_374  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_62 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48_375 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48_375  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_47 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_376 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_376  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [16]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [16]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087 [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0466 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE_377 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE_377  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_DONE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [2]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL_378 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL_378  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0060 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0465 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL_379 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL_379  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0179 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0464 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL_380 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL_380  (
    .I(phyemaccol),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT_381 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT_381  (
    .I(\BU2/U0/N66288 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0463 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED_382 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED_382  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0077 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0462 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_383 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_383  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0076 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0462 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH_384 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH_384  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER_385 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER_385  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0074 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0461 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE_386 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE_386  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0354 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0460 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG_387 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG_387  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0350 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0459 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG_388 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG_388  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0068 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0458 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST_389 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST_389  (
    .I(\BU2/U0/N66185 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0457 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK_390 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK_390  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0456 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH_391 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH_391  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0171 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0455 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD_392 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD_392  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0060 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0454 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD_393 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD_393  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0319 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0453 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH_394 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH_394  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0313 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0452 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS_395 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS_395  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0308 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0451 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_396 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_396  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0167 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0450 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL_397 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL_397  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0302 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0449 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA_398 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA_398  (
    .I(\BU2/U0/N66126 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_399 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_399  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0165 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0448 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_400 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_400  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0296 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0447 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS_401 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS_401  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0291 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0446 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL_402 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL_402  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0287 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0445 ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100_403 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100_403  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0038 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100.GSR.OR ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0001 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7_404 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7_404  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7  (
    .I(clientemactxifgdelay_3[7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN_405 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN_405  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_406 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_406  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0443 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN_407 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN_407  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN_408 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN_408  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE_409 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE_409  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_2 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0063 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [2]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REGPREDELGEN .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REGPREDELGEN  (
    .CLK(txcoreclk),
    .A0(\BU2/U0/address_valid_early ),
    .A1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\BU2/U0/address_valid_early ),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CE(\BU2/U0/address_valid_early ),
    .D(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .Q(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DELAYED ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REGPREDELGEN_Q15_UNCONNECTED )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1_410 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1_410  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt_411 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt_411  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<4>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[9] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<5>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<4>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<3>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<2>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<1>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<0>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN_412 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN_412  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4_413 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4_413  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt_414 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt_414  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<8>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<7>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<6>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6_415 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6_415  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD1 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [6]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [7]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5_416 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5_416  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<2>1 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [29]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<1>1 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [30]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01041 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01041  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0104 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<0>1 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [31]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0063_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0063_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0299 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .O(\BU2/U0/N65592 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER40 .INIT = 16'hAAAB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ER40  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .O(\BU2/U0/CHOICE3268 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00601 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00601  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0060 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01111 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01111  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0111 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0_417 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0_417  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1_418 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1_418  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<5>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<3>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<2>1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<1>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<0>1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<7>1 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<6>1 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<4>1 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2_419 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2_419  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [9]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION_420 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION_420  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0153 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0531 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<13>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<13>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[18] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<1>1 .INIT = 16'hABA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<0>1 .INIT = 16'hABA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<7>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<6>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<5>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<4>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<3>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<2>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<1>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<0>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [5]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [6]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [4]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [5]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [3]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [4]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00681 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00681  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0068 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<7>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<7>1 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [24]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<5>1 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [5]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6_421 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6_421  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01231 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01231  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0123 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<13>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<13>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [13])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt_422 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt_422  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG49 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG49  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [6]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT [7]),
    .O(\BU2/U0/CHOICE2243 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00547 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00547  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [4]),
    .O(\BU2/U0/CHOICE2087 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001146 .INIT = 8'h0E;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n001146  (
    .ADR0(\BU2/U0/CHOICE2209 ),
    .ADR1(\BU2/U0/CHOICE2216 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0011 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125_SW0 .INIT = 16'h7EFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [8]),
    .O(\BU2/U0/N65984 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[25]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<12>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<12>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [12])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<11>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<11>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [11])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<10>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<10>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [10])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<9>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<9>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [9])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<8>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<8>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<7>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<6>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<5>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<4>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<3>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<2>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<1>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<0>1 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00761 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00761  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0076 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_CONTROL1 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_CONTROL1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21490 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [11]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_CONTROL )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<2> .INIT = 16'h8DD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<2>  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [2]),
    .ADR3(\BU2/U0/N51861 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00741 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00741  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0074 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01911 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01911  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0191 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0100<3>1 .INIT = 16'hFF7F;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0100<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21490 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [0]),
    .ADR3(\BU2/U0/N53396 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0100 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01461 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01461  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0146 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3_423 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3_423  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt_424 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt_424  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<0>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4_425 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4_425  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01151 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01151  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0115 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<4>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4374 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<1>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<2>_SW0 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<2>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .O(\BU2/U0/N51861 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<9>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<9>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [9])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<7>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<5>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<4>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<2>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<1>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_391 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_391  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_39 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt_426 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt_426  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC2_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5_427 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5_427  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<3> .INIT = 16'h2772;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<3>  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [3]),
    .ADR3(\BU2/U0/N52182 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01571 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01571  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_ACK_EARLY_IN )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<3>_SW0 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<3>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [1]),
    .O(\BU2/U0/N52182 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01591 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01591  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[1] ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[2] )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [3])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001427 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001427  (
    .ADR0(\BU2/U0/CHOICE2045 ),
    .ADR1(\BU2/U0/CHOICE2048 ),
    .O(\BU2/U0/CHOICE2049 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<5>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[10] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01651 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01651  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0165 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<0>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01671 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01671  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0167 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<1>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG93 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG93  (
    .ADR0(\BU2/U0/CHOICE2243 ),
    .ADR1(\BU2/U0/CHOICE2250 ),
    .ADR2(\BU2/U0/CHOICE2230 ),
    .ADR3(\BU2/U0/CHOICE2237 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED_PRE_REG )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [4]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [4])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n0036_428 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n0036_428  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .ADR1(\BU2/U0/N59033 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_SW14 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_SW14  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [3]),
    .O(\BU2/U0/CHOICE1339 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01741 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01741  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0174 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<2>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<3>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01771 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01771  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0177 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01821 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01821  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01831 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01831  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<4>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [5]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00951 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00951  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0095 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01861 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01861  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0226 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0186 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_431 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_431  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_43 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01881 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01881  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0188 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01891 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01891  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0189 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0063_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0063_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65592 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0063 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01961 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01961  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0196 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01921 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01921  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0192 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<4>1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<5>1 .INIT = 8'hE0;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00111 .INIT = 8'hBF;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n00111  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0011 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_241 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_241  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_24 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<5>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02001 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02001  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0200 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt_429 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt_429  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02021 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02021  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ),
    .ADR2(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0202 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<6>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt_430 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt_430  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<4>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<7>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_68_431  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_67 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_62 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_68 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_45_432  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_45 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_45 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_50_433  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_49 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_45 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_50 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<3>1 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [28]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5_434 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5_434  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>57 .INIT = 16'hE200;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>57  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [10]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19436 ),
    .O(\BU2/U0/CHOICE3012 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_56_435  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_56 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_61 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_56 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2_436 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2_436  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3_437 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3_437  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6_438 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6_438  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5_439 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5_439  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_59_440  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_59 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_64 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_59 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_65_441  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_64 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_59 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_65 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<6>1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01981 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01981  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0198 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_66_442  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_65 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_60 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_66 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_601 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_601  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_60 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<3>1 .INIT = 16'hABA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004540_SW0 .INIT = 16'hEEE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004540_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_N22904 ),
    .ADR2(\BU2/U0/CHOICE2540 ),
    .ADR3(\BU2/U0/CHOICE3280 ),
    .O(\BU2/U0/N65759 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_611 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_611  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_61 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_60_443  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_60 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_65 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_60 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0  (
    .I(clientemactxifgdelay_3[0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [2]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [2]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_631 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_631  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_63 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_62_444  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_62 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_67 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_62 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt_445 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt_445  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2  (
    .I(clientemactxifgdelay_3[2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3  (
    .I(clientemactxifgdelay_3[3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6_446 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6_446  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_49_447  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_48 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_44 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_49 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6  (
    .I(clientemactxifgdelay_3[6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_DONE1 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_DONE1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_DONE )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n025614_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n025614_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [5]),
    .O(\BU2/U0/N65420 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02571 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02571  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_441 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_441  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_45 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_44 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49_448 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49_448  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_48 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087 [0]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [0]),
    .CE(VCC),
    .RST(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_48_449  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_48 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<4>1 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_OUT<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0026 [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [27]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0_450 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0_450  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_461 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_461  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_46 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012171 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012171  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN__n0108 [1]),
    .ADR1(\BU2/U0/CHOICE2940 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN__n0106 [1]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0012 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_46_451  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_46 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_46 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2_452 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2_452  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1_453 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1_453  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1 ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_51_454  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_50 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_46 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_51 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12_455 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12_455  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13_456 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13_456  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02731 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02731  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0273 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_471 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_471  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_47 )
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11_457 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11_457  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n031923 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n031923  (
    .ADR0(\BU2/U0/CHOICE2424 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [0]),
    .ADR3(\BU2/U0/CHOICE2430 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0319 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_52_458  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_51 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_47 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_52 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [1]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [0]),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_641 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_641  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_64 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_53_459  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_52 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_48 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_53 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_481 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_481  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_48 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4_460 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4_460  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_47_461  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_47 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_51 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_47 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53_462 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53_462  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_52 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_53 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_491 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_491  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_49 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_48_463  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_48 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_52 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_48 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54_464 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54_464  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_53 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [6]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_49_465  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_49 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_53 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_49 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11_466 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11_466  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148856_SW1 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker2148856_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [10]),
    .O(\BU2/U0/N65882 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55_467 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55_467  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_54 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[2] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56_468 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56_468  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_55 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_56 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04491 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04491  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0302 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0449 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_45_469 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_45_469  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_44 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_45 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03021 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03021  (
    .ADR0(\BU2/U0/TRIMAC_INST_INT_TX_UNDERRUN_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR2(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0302 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57_470 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57_470  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_56 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58_471 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58_471  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_57 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_58 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<12>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<12>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[17] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6_472 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6_472  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03081 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03081  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21290 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0308 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59_473 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59_473  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_58 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<11>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<11>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[16] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47_474 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47_474  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_46 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_46_475 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_46_475  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_45 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_46 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60_476 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60_476  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_59 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03151 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n03151  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0315 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65_477 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65_477  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_64 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64_478 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64_478  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_63 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_64 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001426 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001426  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [8]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [9]),
    .O(\BU2/U0/CHOICE2048 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61_479 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61_479  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_60 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_61 ),
    .SET(GND),
    .RST(GSR)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_56_480  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_55 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_50 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_56 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt_481 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt_481  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q1_ASSIGN_LI_rt ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_55_482  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/N66317 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_55 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt_483 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt_483  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC5_Q<0>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<10>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<10>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[15] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62_484 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62_484  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_61 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_62 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<8>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<8>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[13] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_50_485  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_50 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_55 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_50 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0_486 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0_486  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6_487 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6_487  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5_488 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5_488  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0113 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<9>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<9>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[14] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9_489 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9_489  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2_490 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2_490  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN__n003331 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN__n003331  (
    .ADR0(\BU2/U0/CHOICE2117 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6 [4]),
    .ADR3(\BU2/U0/N65452 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN__n0033 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0_491 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0_491  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[12] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1_492 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1_492  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1 ),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_51_493  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_51 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_56 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_51 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_57_494  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_56 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_51 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_57 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<6>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[11] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2_495 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2_495  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_59_496  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_58 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_53 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_59 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_52_497  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_52 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_57 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_52 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_58_498  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_57 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_52 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_58 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3_499 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3_499  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [3]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_53_500  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_53 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_58 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_53 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001290 .INIT = 16'hFF90;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO__n001290  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .ADR3(\BU2/U0/CHOICE3181 ),
    .O(\BU2/U0/CHOICE3182 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4_501 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4_501  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [5]),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_60_502  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_59 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_54 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_60 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1_503 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1_503  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_54_504  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_54 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_59 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_54 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4_505 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4_505  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_55 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5_506 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5_506  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_61_507  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_60 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_55 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_61 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3_508 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3_508  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_54 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6_509 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6_509  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6 ),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_55_510  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_55 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_60 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_55 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00771 .INIT = 16'h00AE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00771  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0177 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0077 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7_511 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7_511  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8_512 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8_512  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<4>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9_513 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9_513  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<6>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3_514 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3_514  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3 ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_62_515  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_61 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_56 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_62 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<5>1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0040_Result<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0161 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0040 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10_516 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10_516  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<2>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<3>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2  (
    .I(\BU2/U0/address_valid_early ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST [2]),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_63_517  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_62 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_57 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_63 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE [13]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12_518 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12_518  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12 ),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_57_519  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_57 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_62 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_57 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<18>1 .INIT = 16'hD888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<18>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [9]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [18]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [18])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4_520 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4_520  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02877 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n02877  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE ),
    .O(\BU2/U0/CHOICE2778 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13_521 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13_521  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4370 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_ClkEn_INV1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_ClkEn_INV1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0_522 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0_522  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_64_523  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_63 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_58 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_64 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<8>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<8>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1_524 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1_524  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<0>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[5] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2_525 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2_525  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_591 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_591  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_59 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_58_526  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_58 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_63 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_58 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<1>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[6] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3_527 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3_527  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0112 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0_528 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0_528  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0114 [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[7] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4_529 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4_529  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5_530 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5_530  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1  (
    .I(clientemactxifgdelay_3[1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6_531 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6_531  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6 ),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_67_532  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_66 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_61 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_67 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux_INT_BYTE_COUNT_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[8] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7_533 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7_533  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8_534 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8_534  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [8]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9_535 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9_535  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [9]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10_536 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10_536  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [10]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11_537 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11_537  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [11]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12_538 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12_538  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [12]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_621 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_621  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .ADR1(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_63 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_62 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_61_539  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_61 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_66 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_61 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00841 .INIT = 16'h888A;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n00841  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0218 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13_540 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13_540  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0134 [13]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_N5803 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8_541 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8_541  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_59 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04271 .INIT = 8'h07;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04271  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0427 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0_542 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0_542  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_51 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01531 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n01531  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0153 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1_543 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1_543  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_52 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1 ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4  (
    .I(clientemactxifgdelay_3[4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3_544 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3_544  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3 ),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_63_545  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_63 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_68 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_sum_63 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_69_546  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_68 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_lut3_63 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_inst_cy_69 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50_547 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50_547  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_49 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0468 ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_44_548  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_44 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_cy_48 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_sum_44 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_451 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_451  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0386 ),
    .ADR1(\BU2/U0/address_valid_early ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_46 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_inst_lut3_45 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04431 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04431  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0443 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<2>1 .INIT = 16'hC9FF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<1>1 .INIT = 8'hD7;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<0>1 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0083 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029118 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n029118  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ),
    .O(\BU2/U0/CHOICE3129 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087<1>1 .INIT = 8'hD7;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087<0>1 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0087 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088<1>1 .INIT = 8'hD7;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088<0>1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0088 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00451 .INIT = 16'hABAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00451  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ),
    .ADR2(\BU2/U0/CHOICE1339 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<11>161_G .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<11>161_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [5]),
    .O(\BU2/U0/N66084 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025_549 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025_549  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .ADR1(\BU2/U0/N50430 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04501 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04501  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0167 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0450 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04511 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04511  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0308 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0451 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04521 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04521  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0313 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0452 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00541 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00541  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .ADR2(\BU2/U0/CHOICE2257 ),
    .ADR3(\BU2/U0/CHOICE2262 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0054 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000874 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000874  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ),
    .O(\BU2/U0/CHOICE2709 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025_SW0 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0025_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD ),
    .O(\BU2/U0/N50430 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04561 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04561  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0315 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0336 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0456 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04571 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04571  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0173 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0457 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0158 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0158  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH ),
    .ADR3(\BU2/U0/N51266 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[1] )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010212_G .INIT = 16'hF200;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0010212_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Msub__n0022__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_OCCUPANCY [1]),
    .ADR2(\BU2/U0/CHOICE3286 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .O(\BU2/U0/N66089 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04641 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04641  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR1(\BU2/U0/N65254 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DELAYED ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0464 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00052 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00052  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [6]),
    .O(\BU2/U0/CHOICE3329 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05311 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05311  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0531 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04671 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04671  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_TIME_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0467 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014_SW0 .INIT = 16'hFEFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0014_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME ),
    .O(\BU2/U0/N50821 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16_SW1 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .O(\BU2/U0/N65478 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<17>1 .INIT = 16'hD888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<17>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [17]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [17])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<16>1 .INIT = 16'hD888;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<16>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [16]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [16])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0158_SW0 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0158_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH ),
    .O(\BU2/U0/N51266 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt_550 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt_550  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [8]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_LENGTH_CNT<8>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_3 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0062 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [3]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04701 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04701  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_65 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21500 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0470 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04711 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04711  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_60 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0471 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04721 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04721  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_COUNT_57 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0472 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04731 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04731  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0226 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0256 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0273 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0473 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04741 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04741  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0474 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046173_SW0 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n046173_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/N65408 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05101 .INIT = 16'hFF2F;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05101  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_BURSTING ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0510 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_STATUS_VECTOR[1] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<10>161_G .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<10>161_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [4]),
    .O(\BU2/U0/N66094 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05141 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05141  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0514 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[7] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05131 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05131  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21525 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR2(\BU2/U0/TRIMAC_INST_INT_TX_UNDERRUN_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0513 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00211 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00211  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0021 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[26]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05231 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05231  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0523 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05241 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05241  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_EXCESSIVE_COLLISIONS ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0524 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05251 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05251  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0525 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<16>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED<7>_rt1 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0538<15>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[16] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4600 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0215<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0215 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0039 [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt_551 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt_551  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05271 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05271  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0527 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05281 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05281  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0528 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[27]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<18>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4538 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0224<17>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [18])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05301 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05301  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0530 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06721 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06721  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [3]),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06731 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06731  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [2]),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06741 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06741  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [1]),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN_552 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN_552  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stagecy_rn_6  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Eq_stage_cyo6 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4625 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0226 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06751 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n06751  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_RETRY [0]),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_4 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0061 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [4]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<14>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N4442 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0245<13>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0245 [14])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[28]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010_553 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010_553  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0022 ),
    .ADR2(\BU2/U0/N52675 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Ker21493  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1 ),
    .ADR3(\BU2/U0/N51500 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_N21495 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<0>16 .INIT = 8'h72;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<0>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010_SW0 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n0010_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7 ),
    .O(\BU2/U0/N52675 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<8>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<8>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<7>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<6>1 .INIT = 16'hFFB8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [4])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<9>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT<9>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_STATE_MACH__n0246<8>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [9])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5  (
    .I(clientemactxifgdelay_3[5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1__n0000 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[0] ),
    .CE(VCC),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mxor__n0000_Result1 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mxor__n0000_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[14] ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00471 .INIT = 16'h2AAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00471  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [0]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>162 .INIT = 16'h01D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_Mmux_WR_OCCUPANCY_Result<2>162  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .O(\BU2/U0/CHOICE1804 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Ker171201 .INIT = 4'h7;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Ker171201  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_47 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_N17122 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00491 .INIT = 16'hA2AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00491  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_N17122 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[14] ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [2]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [3]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [4]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [5]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [6]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [7]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29_554 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29_554  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>__net3 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29 ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00331 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00331  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_N17122 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [9])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00351 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00351  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [1]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00391 .INIT = 16'h222A;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00391  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [6]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_48 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [6])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00411 .INIT = 16'h22A2;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00411  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_N17122 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00431 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC__n00431  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_50 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ATTEMPT_COUNT_49 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_srl_0 .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_srl_0  (
    .CLK(txcoreclk),
    .A0(\BU2/U0/address_valid_early ),
    .A1(\BU2/U0/address_valid_early ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A3(\BU2/U0/address_valid_early ),
    .CE(\BU2/U0/address_valid_early ),
    .D(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[0] ),
    .Q(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>__net3 ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_srl_0_Q15_UNCONNECTED )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0059_Result_SW1 .INIT = 16'h9669;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0059_Result_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0296 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0295 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [26]),
    .O(\BU2/U0/N65768 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [8]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q [0]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TC ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TC ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TC ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [1]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I291  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C7 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ7 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I278  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<6>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C6 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ6 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I265  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<5>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C5 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ5 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I252  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<4>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C4 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ4 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I239  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<3>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ3 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I226  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<2>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C2 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ2 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<1>_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ1 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_C7 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TC )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I250 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I250 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I250  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ4 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [4]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I224 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I224 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I224  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ2 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [2]),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TC ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I289 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I289 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I289  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ7 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q7_ASSIGN_LI ),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I276 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I276 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I276  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ6 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [6]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I263 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I263 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I263  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ5 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [5]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I36 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [0]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I35 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I35  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ1 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF6  (
    .I(\BU2/U0/address_valid_early ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6q ),
    .SET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5q ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TC_ASSIGN_I0 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int6 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I36  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TQ0 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI ),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_Q0_ASSIGN_LI_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_TQ0 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5q ),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I298  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_C1 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TC )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC4_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int3q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC3_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int2q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC2_Q [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_FF1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1 ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int1q ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I237 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I237 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_X36_1I237  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_TQ3 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE ),
    .RST(GSR),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [3]),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I6  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ0 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I28  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_Q1_ASSIGN_LI_rt ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_C1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TQ1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_24_555  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_24 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_26 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_24 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_27_556  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_26 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_24 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_27 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_23_557  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_23 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_25 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_23 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_26_558  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_25 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_23 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_26 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_22_559  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_22 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_24 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_22 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_25_560  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_24 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_22 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_25 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_24_561  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/N66312 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_24 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_25_562  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_25 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_27 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_25 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [2]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [3]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_281 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_281  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_RD_ADV ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[5] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_28 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_30_563  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_29 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_27 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_30 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [1]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [2]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt_564 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt_564  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<3>_rt ),
    .ADR1(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_29_565  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_28 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_26 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_29 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN<5>1 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN<5>1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(corehassgmii),
    .ADR2(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[5] )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000057_SW1 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n000057_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [9]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [10]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [12]),
    .O(\BU2/U0/N65878 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR [0]),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [1]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_26 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_26 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_26  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_26 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [4])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_25 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_25 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_25  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_25 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [3])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_23 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_23  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_23 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [1])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_22 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_22  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_22 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN<3>1 .INIT = 8'hBF;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN<3>1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(corehassgmii),
    .ADR2(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_DIN[3] )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_26_566  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_26 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_28 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_26 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_28_567  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_28 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_30 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_28 )
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_28 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_28 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_28  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_28 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [6])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_27 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_27 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_27  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_27 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [5])
  );
  initial assign \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_24 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_24 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_24  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_24 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(GSR),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT [2])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_27_568  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_27 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_29 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_sum_27 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_4  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [4]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [4]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_3  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [3]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [3]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_2  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [2]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [2]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [1]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [0]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_10  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [10]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [10]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N48701 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N48701  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2_569 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2_569  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1_570 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1_570  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In46 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In46  (
    .ADR0(\BU2/U0/CHOICE2384 ),
    .ADR1(\BU2/U0/N65472 ),
    .ADR2(\BU2/U0/CHOICE2389 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt_571 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt_571  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC1_Q<3>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<8>_SW0 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<8>_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[17] ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0538[8] ),
    .O(\BU2/U0/N56896 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_11  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [11]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [11]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<12>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<12>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [12]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4156 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4152 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [11])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4152 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [11]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4152 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4148 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [10])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4148 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<10>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [10]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4148 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4144 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [9])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4144 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<9>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [9]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4144 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4140 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [8])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4140 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<8>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4140 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4136 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [7])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4136 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [7]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4136 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4132 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [6])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4132 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<6>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [6]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4132 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4128 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [5])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4128 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<5>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [5]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4128 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4124 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [4])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4124 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<4>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [4]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4124 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4120 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [3])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4120 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<3>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4120 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4116 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4116 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<2>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [2]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4116 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4112 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [1])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4112 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<1>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [1]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4112 ),
    .ADR1(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt ),
    .I1(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [0])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>cy  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER<0>_rt ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<0>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_6  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [6]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [6]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_Ker127001 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_Ker127001  (
    .ADR0(\BU2/U0/N66330 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N12702 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_7  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [7]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [7]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<8> .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_Mmux__n0001_Result<8>  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0084 ),
    .ADR1(\BU2/U0/N56896 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0002 [8]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT__n0001 [8])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_12  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [12]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [12]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_572 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_572  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0004 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING ),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3_573 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3_573  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3-In ),
    .SET(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_9  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [9]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [9]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_8  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [8]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [8]),
    .SET(GND),
    .RST(GSR)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<12>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_N4156 ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_BURST_STATE_MACH__n0006<11>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0006 [12])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<0>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<0>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [8]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT_574 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT_574  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0012 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT_575 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT_575  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0011 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0__n00011 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0001 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_28_576  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_27 ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_lut3_25 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_RATE_GEN_COUNT_inst_cy_28 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_BYTECNTSRL .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_TXGEN_BYTECNTSRL  (
    .CLK(txcoreclk),
    .A0(\BU2/U0/address_valid_early ),
    .A1(\BU2/U0/address_valid_early ),
    .A2(\BU2/U0/address_valid_early ),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CE(\BU2/U0/address_valid_early ),
    .D(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .Q(\BU2/U0/TRIMAC_INST_TXGEN_INT_TX_EN_DELAY ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_TXGEN_BYTECNTSRL_Q15_UNCONNECTED )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA_14  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_Mshreg_SHIFT_DATA<13>_29 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_prbs_1_SHIFT_DATA[14] ),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0005 [5]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_INT_BURSTING_N4870 ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_BURST_COUNTER [5]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4_577 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4_577  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4-In ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_5 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG_5  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0060 ),
    .SRST(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_REG [5]),
    .SET(GND),
    .RST(GSR),
    .SSET(GND)
  );
  X_AND2 \BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_X36_1I956  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int4q ),
    .I1(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_CRC5_TC ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRCGEN2_int5 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN_578 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN_578  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0016 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT_579 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT_579  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0017 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT_580 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT_580  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0018 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT_581 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT_581  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0019 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT_582 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT_582  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0020 ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT_583 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT_583  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT_584 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT_584  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0013 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT_585 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT_585  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0014 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRC_CE1 .INIT = 16'hB8BB;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_CRC_CE1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN ),
    .ADR1(tieemacconfigvec_7[66]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN ),
    .ADR3(tieemacconfigvec_7[65]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRC_CE )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [1]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT_586 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT_586  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG_587 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG_587  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR [0]),
    .CE(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES_PRE_REG1 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES_PRE_REG1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_INT_TX_EN_DELAY ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES_PRE_REG )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00111 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN__n00111  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0011 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00121 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00121  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<1>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<1>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [9]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00141 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00141  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<4>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<4>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [12]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00161 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN__n00161  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0016 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00171 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN__n00171  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0017 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00181 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00181  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0018 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<2>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [10]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00201 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00201  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0020 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN_588 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN_588  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0022 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_CRS_589 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_CRS_589  (
    .I(phyemaccrs),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE_590 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE_590  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN__n0034 ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<3>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [11]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00221 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN__n00221  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0022 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00131 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00131  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0013 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX_591 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX_591  (
    .I(tieemacconfigvec_7[55]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100_592 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100_592  (
    .I(NlwRenamedSig_OI_speedis10100),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE_593 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE_593  (
    .I(tieemacconfigvec_7[59]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE_594 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE_594  (
    .I(tieemacconfigvec_7[57]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE_595 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE_595  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_VLAN_ENABLE_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN_596 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN_596  (
    .I(tieemacconfigvec_7[54]),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES_PRE_REG ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[30]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<7>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [15]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TX_EN_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TX_EN_Result1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [1]),
    .O(\BU2/U0/TRIMAC_INST__n0011 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG_597 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG_597  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT ),
    .RST(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00191 .INIT = 8'h8A;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN__n00191  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0019 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<5>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<5>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [13]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TX_ER_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TX_ER_Result1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [1]),
    .O(\BU2/U0/TRIMAC_INST__n0012 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_EXTENSION_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_EXTENSION_Result1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0039 [1]),
    .O(\BU2/U0/TRIMAC_INST_INT_EXTENSION )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN__n00341 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN__n00341  (
    .ADR0(tieemacconfigvec_7[58]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN__n0034 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<6>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_Mmux_TXD_Result<6>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [14]),
    .O(\BU2/U0/TRIMAC_INST__n0009 [6])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<1>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [1]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [1])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<0>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [0]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [0])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [6]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [5]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [4]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [3]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [2]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [1]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<3>1 .INIT = 8'h06;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n0007 [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX__n0012 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [3])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<2>1 .INIT = 16'h006A;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX__n0012 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<1>1 .INIT = 8'h06;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX__n0012 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>0 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<9>0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q [0]),
    .O(\BU2/U0/CHOICE1945 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14  (
    .I(clientemacpauseval_4[14]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13  (
    .I(clientemacpauseval_4[13]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12  (
    .I(clientemacpauseval_4[12]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11  (
    .I(clientemacpauseval_4[11]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10  (
    .I(clientemacpauseval_4[10]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9  (
    .I(clientemacpauseval_4[9]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8  (
    .I(clientemacpauseval_4[8]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7  (
    .I(clientemacpauseval_4[7]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6  (
    .I(clientemacpauseval_4[6]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5  (
    .I(clientemacpauseval_4[5]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4  (
    .I(clientemacpauseval_4[4]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3  (
    .I(clientemacpauseval_4[3]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2  (
    .I(clientemacpauseval_4[2]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1  (
    .I(clientemacpauseval_4[1]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0  (
    .I(clientemacpauseval_4[0]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2_598 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2_598  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1_599 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1_599  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1-In ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt_600 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt_600  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q [6]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC3_Q<6>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In30 .INIT = 16'hFFE0;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In30  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR1(\BU2/U0/CHOICE2173 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .ADR3(\BU2/U0/CHOICE2177 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2-In )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<3>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [11]),
    .O(\BU2/U0/CHOICE2833 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [4]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25  (
    .I(tieemacconfigvec_7[25]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [25]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28  (
    .I(tieemacconfigvec_7[28]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [28]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27  (
    .I(tieemacconfigvec_7[27]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [27]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30  (
    .I(tieemacconfigvec_7[30]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [30]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29  (
    .I(tieemacconfigvec_7[29]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [29]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15  (
    .I(tieemacconfigvec_7[15]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14  (
    .I(tieemacconfigvec_7[14]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23  (
    .I(tieemacconfigvec_7[23]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [23]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22  (
    .I(tieemacconfigvec_7[22]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [22]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21  (
    .I(tieemacconfigvec_7[21]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [21]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31  (
    .I(tieemacconfigvec_7[31]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [31]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n00011 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n00011  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n0007 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6  (
    .I(tieemacconfigvec_7[6]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24  (
    .I(tieemacconfigvec_7[24]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [24]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46  (
    .I(tieemacconfigvec_7[46]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [46]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<4>1 .INIT = 16'h006A;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Madd__n0000__n0007 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX__n0012 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [4])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26  (
    .I(tieemacconfigvec_7[26]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [26]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG_601 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG_601  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0066 ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3_602 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3_602  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3-In ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .CE(VCC),
    .RST(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_ACK_OUT2  (
    .IA(\BU2/U0/TRIMAC_INST_INT_TX_ACK_EARLY_IN ),
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .O(\NLW_BU2/U0/TRIMAC_INST_FLOW_TX_MUX_ACK_OUT2_O_UNCONNECTED )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_ACK_OUT  (
    .IA(\BU2/U0/TRIMAC_INST_INT_TX_ACK_IN ),
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_COMB )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_CONTROL_COMPLETE1 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_CONTROL_COMPLETE1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_CONTROL_COMPLETE )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT_603 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT_603  (
    .I(\BU2/U0/TRIMAC_INST_INT_TX_ACK_IN ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47  (
    .I(tieemacconfigvec_7[47]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [47]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<0>1 .INIT = 8'h01;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR2(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11  (
    .I(tieemacconfigvec_7[11]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194161 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194161  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19418 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<6>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [38]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_N19412 ),
    .ADR2(\BU2/U0/N66190 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [46]),
    .O(\BU2/U0/CHOICE3091 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00057 .INIT = 16'h8000;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN__n00057  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [3]),
    .O(\BU2/U0/CHOICE3332 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125_SW1 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<0>125_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [24]),
    .O(\BU2/U0/N65986 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000857 .INIT = 16'hF200;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER__n000857  (
    .ADR0(\BU2/U0/CHOICE2702 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD ),
    .ADR2(\BU2/U0/CHOICE2693 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA ),
    .O(\BU2/U0/CHOICE2706 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>4 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<2>4  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [34]),
    .ADR1(\BU2/U0/N66135 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [42]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_N19406 ),
    .O(\BU2/U0/CHOICE2998 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00544 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00544  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [5]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .O(\BU2/U0/CHOICE2085 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD_604 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD_604  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0067 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5  (
    .I(tieemacconfigvec_7[5]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00241 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00241  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ),
    .ADR3(\BU2/U0/CHOICE1339 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0024 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4  (
    .I(tieemacconfigvec_7[4]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00221 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n00221  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0022 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n045423 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n045423  (
    .ADR0(\BU2/U0/N66248 ),
    .ADR1(\BU2/U0/CHOICE2651 ),
    .ADR2(\BU2/U0/CHOICE2655 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0454 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1  (
    .I(tieemacconfigvec_7[1]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0  (
    .I(tieemacconfigvec_7[0]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7  (
    .I(tieemacconfigvec_7[7]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2  (
    .I(tieemacconfigvec_7[2]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8  (
    .I(tieemacconfigvec_7[8]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3  (
    .I(tieemacconfigvec_7[3]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9  (
    .I(tieemacconfigvec_7[9]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10  (
    .I(tieemacconfigvec_7[10]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41  (
    .I(tieemacconfigvec_7[41]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [41]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40  (
    .I(tieemacconfigvec_7[40]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [40]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39  (
    .I(tieemacconfigvec_7[39]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [39]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42  (
    .I(tieemacconfigvec_7[42]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [42]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12  (
    .I(tieemacconfigvec_7[12]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34  (
    .I(tieemacconfigvec_7[34]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [34]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17  (
    .I(tieemacconfigvec_7[17]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [17]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36  (
    .I(tieemacconfigvec_7[36]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [36]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16  (
    .I(tieemacconfigvec_7[16]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [16]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20  (
    .I(tieemacconfigvec_7[20]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [20]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35  (
    .I(tieemacconfigvec_7[35]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [35]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00465 .INIT = 16'hEAAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX__n00465  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .O(\BU2/U0/CHOICE1379 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43  (
    .I(tieemacconfigvec_7[43]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [43]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18  (
    .I(tieemacconfigvec_7[18]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [18]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44  (
    .I(tieemacconfigvec_7[44]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [44]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37  (
    .I(tieemacconfigvec_7[37]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [37]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In_605 .INIT = 16'h00AE;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In_605  (
    .ADR0(\BU2/U0/N60912 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13  (
    .I(tieemacconfigvec_7[13]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38  (
    .I(tieemacconfigvec_7[38]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [38]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19  (
    .I(tieemacconfigvec_7[19]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [19]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45  (
    .I(tieemacconfigvec_7[45]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [45]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32  (
    .I(tieemacconfigvec_7[32]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [32]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15  (
    .I(clientemacpauseval_4[15]),
    .CE(clientemacpausereq),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT_606 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT_606  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0011 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0069 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_COMB ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxack),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021812 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n021812  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [7]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT [4]),
    .O(\BU2/U0/CHOICE2949 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0014 [7]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00041 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX__n00041  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33  (
    .I(tieemacconfigvec_7[33]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX__n0004 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [33]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_607 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_607  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0046 ),
    .CE(\BU2/U0/N66297 ),
    .SET(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<1>1 .INIT = 16'h99F9;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00671 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX__n00671  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .ADR1(\BU2/U0/N66180 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0067 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<7>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [7]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [7])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL_608 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL_608  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX__n0015 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n00691 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n00691  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_CONTROL_COMPLETE ),
    .ADR1(clientemacpausereq),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX__n0069 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194401 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_Ker194401  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_N19442 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG_609 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG_609  (
    .I(clientemactxdvld),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1 .INIT = 16'h2300;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_Mmux__n0001_Result<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [5])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_OUT1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_OUT1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL ),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_UNDERRUN_OUT )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [7]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [7])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<6>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<6>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [6]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [6])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_Ker185151 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_Ker185151  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [4]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_N18517 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0011 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0010 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0009 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0008 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0007 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0014 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0013 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0012 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0011 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0010 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0009 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0008 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0007 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT_610 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT_610  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0004 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0039 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT_611 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT_611  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0004 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0038 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In_612 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In_612  (
    .ADR0(\BU2/U0/N52009 ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3__n0000 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE1 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE1  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME ),
    .O(emacclientrxstats_6[24])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ1 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_PAUSE_REQ_LOCAL )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [4]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00001 .INIT = 16'h0002;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_N18510 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00041 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_RX__n00041  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0004 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00071 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00071  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [7]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0007 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00081 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00081  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [6]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0008 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00091 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00091  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [5]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0009 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00101 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00101  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [4]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0010 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00111 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00111  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [3]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0011 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00121 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00121  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [2]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00131 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00131  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [1]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0013 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00141 .INIT = 8'h10;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX__n00141  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_DATA [0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<1>1 .INIT = 16'h0006;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR2(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR3(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_OUT1 .INIT = 16'hA2AA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_OUT1  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_COMB )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE44 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_DONE44  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [12]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT [11]),
    .O(\BU2/U0/CHOICE2463 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>16 .INIT = 16'h00D8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [1]),
    .ADR3(tieemacconfigvec_7[66]),
    .O(\BU2/U0/CHOICE2325 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<2>1 .INIT = 16'h006A;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01621 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n01621  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0162 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [1]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [1]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_Ker185081 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX_Ker185081  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_N18510 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [2]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [2]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [3]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [3]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [4]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [4]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [5]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [5]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0036 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [0]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [0]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_Ker184871 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_RX_Ker184871  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n0036_SW0 .INIT = 16'hFBFF;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n0036_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [4]),
    .O(\BU2/U0/N59033 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0012 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0013 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX__n0014 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [7]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [7]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00381 .INIT = 16'hEAAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n00381  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_N18510 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX__n0021 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0038 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [6]),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_RX__n0000 ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_OPCODE_EARLY [6]),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00391 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n00391  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_N18489 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_N18510 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX__n0021 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0039 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00491 .INIT = 16'hFEEE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n00491  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR1(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_N18517 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0049 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005129 .INIT = 16'hF888;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n005129  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .ADR2(\BU2/U0/CHOICE2197 ),
    .ADR3(\BU2/U0/CHOICE2201 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0051 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_6 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [6])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_21_613  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_21 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_22 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_21 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17_614 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17_614  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_17 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_211 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_211  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [15]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_21 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_20_615  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_20 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_21 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_20 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_22_616  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_21 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_20 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_22 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_201 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_201  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [14]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_20 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_19_617  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_19 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_20 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_19 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_21_618  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_20 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_19 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_21 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_191 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_191  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [13]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_19 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_18_619  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_18 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_19 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_18 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_20_620  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_19 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_18 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_20 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_181 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_181  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [12]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_18 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_17_621  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_17 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_18 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_17 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_19_622  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_18 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_17 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_19 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_171 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_171  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [11]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_17 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_16_623  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_16 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_17 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_16 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_18_624  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_17 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_16 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_18 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_161 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_161  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [10]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_16 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_15_625  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_15 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_16 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_15 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_17_626  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_16 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_15 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_17 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_151 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_151  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [9]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [15]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_15 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_14_627  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_14 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_15 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_14 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_16_628  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_15 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_14 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_16 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_141 .INIT = 8'h27;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_141  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [8]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [14]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_14 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_13_629  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_13 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_14 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_13 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_15_630  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_14 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_13 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_15 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_12_631  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_12 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_13 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_12 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_14_632  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_13 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_12 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_14 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_11_633  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_11 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_12 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_11 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_13_634  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_12 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_11 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_13 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_10_635  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_10 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_11 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_10 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_12_636  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_11 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_10 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_12 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_9_637  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_9 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_10 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_9 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_11_638  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_10 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_9 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_11 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_8_639  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_8 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_9 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_8 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_10_640  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_9 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_8 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_10 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_7_641  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_7 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_8 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_7 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_9_642  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_8 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_7 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_9 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_6_643  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_6 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_7 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_6 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_8_644  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_7 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_lut3_6 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_8 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_7_645  (
    .IB(\BU2/U0/address_valid_early ),
    .SEL(\BU2/U0/N66116 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_cy_7 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21_646 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21_646  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_21 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20_647 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20_647  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_20 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_3 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [3])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_2 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [2])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_1 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [1])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_0 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_5_648  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_5 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_5 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_5 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18_649 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18_649  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_18 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_421 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_421  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_42 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_4_650  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_4 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_4 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_4 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_5_651  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_4 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_4 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_5 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_411 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_411  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_41 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_3_652  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_3 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_3 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_4_653  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_3 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_3 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_4 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_401 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_401  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_40 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_2_654  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_2 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_2 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_2 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_3_655  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_2 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_2 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_3 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<0>1 .INIT = 16'h00A8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [0])
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_1_656  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_1 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_1 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_1 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_2_657  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_1 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_1 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_2 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_381 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_381  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_38 )
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_0_658  (
    .I0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_0 ),
    .I1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_0 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_0 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_1_659  (
    .IB(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_0 ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_lut3_0 ),
    .IA(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_1 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_371 .INIT = 8'h2A;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_371  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_inst_lut3_37 )
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_0_660  (
    .IB(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SEL(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0008 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_cy_0 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<4>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<4>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [4]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [4])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_5 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [5])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<0>1 .INIT = 8'h07;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT ),
    .ADR1(\BU2/U0/CHOICE2600 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00081 .INIT = 4'h8;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00081  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0008 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_13 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [13])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_12 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [12])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG_661 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG_661  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001162 .INIT = 16'h0001;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001162  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20 ),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21 ),
    .O(\BU2/U0/CHOICE2501 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_9 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [9])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001447 .INIT = 16'hAAA8;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001447  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0002 ),
    .ADR1(\BU2/U0/CHOICE2038 ),
    .ADR2(\BU2/U0/CHOICE2041 ),
    .ADR3(\BU2/U0/CHOICE2049 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0014 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_10 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [10])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_14 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [14])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_15 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [15])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_11 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [11])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16_662 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16_662  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_16 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In_SW0 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2-In_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3 ),
    .ADR1(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/N60912 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW__n00071 .INIT = 16'hAEAA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW__n00071  (
    .ADR0(NlwRenamedSig_OI_emacclienttxstatsvld),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [0]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [1]),
    .O(\BU2/U0/TRIMAC_INST_FLOW__n0007 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00221 .INIT = 8'hEA;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n00221  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0011 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0022 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19_663 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19_663  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_19 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_664 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_664  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0014 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0021 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG_665 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG_665  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG ),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_666 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_666 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_666  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_8 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [8])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT_667 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT_667  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0007 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0022 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_inst_sum_4 ),
    .CE(\BU2/U0/address_valid_early ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA [4])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [13]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [13]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [12]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [12]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [11]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [11]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [10]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [10]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [9]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [9]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [8]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [8]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [7]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [7]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [6]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [6]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [5]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [5]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [4]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [4]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [3]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [2]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [1]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [0]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX_668 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX_668  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_PAUSE_REQ_LOCAL ),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [15]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [15]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX_669 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX_669  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE__n0000 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3_670 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3_670  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2_671 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2_671  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1_672 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1_672  (
    .I(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE__n00001 .INIT = 8'hFE;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE__n00001  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3 ),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE__n0000 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [4]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [3]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [2]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [1]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6  (
    .I(clientemactxd_2[6]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5  (
    .I(clientemactxd_2[5]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4  (
    .I(clientemactxd_2[4]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3  (
    .I(clientemactxd_2[3]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2  (
    .I(clientemactxd_2[2]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1  (
    .I(clientemactxd_2[1]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0  (
    .I(clientemactxd_2[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_COMB ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxbadframe),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_COMB ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxgoodframe),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxdvld),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [7]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_inst_sum_7 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n0020 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT [7])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14  (
    .I(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE [14]),
    .CE(NlwRenamedSig_OI_emacclientrxstats[0]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [14]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<5>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<5>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [5]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [5])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In_SW0 .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1-In_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER ),
    .O(\BU2/U0/N52009 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7  (
    .I(clientemactxd_2[7]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [7]),
    .CE(VCC),
    .SET(GND)
  );
  X_XOR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<2>_xor  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4358 ),
    .I1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<1>_cyo ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0004 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_VLAN_ENABLE_OUT1 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW_TX_VLAN_ENABLE_OUT1  (
    .ADR0(tieemacconfigvec_7[56]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_VLAN_ENABLE_OUT )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW__n00011 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW__n00011  (
    .ADR0(NlwRenamedSig_OI_emacclienttxstatsvld),
    .O(\BU2/U0/TRIMAC_INST_FLOW__n0001 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW__n00021 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW__n00021  (
    .ADR0(tieemacconfigvec_7[62]),
    .ADR1(tieemacconfigvec_7[48]),
    .O(\BU2/U0/TRIMAC_INST_FLOW__n0002 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW__n00031 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_FLOW__n00031  (
    .ADR0(tieemacconfigvec_7[61]),
    .ADR1(tieemacconfigvec_7[55]),
    .O(\BU2/U0/TRIMAC_INST_FLOW__n0003 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [5]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [3]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [3])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00591 .INIT = 16'hFF2F;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n00591  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6 ),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM__n0059 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT_673 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT_673  (
    .I(clientemactxunderrun),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<5>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<5>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [5]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [5]),
    .O(emacphytxd_0[5])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_DATA [6]),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6.GSR.OR ),
    .CLK(rxcoreclk),
    .O(emacclientrxd_5[6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxretransmit),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT  (
    .I(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxcollision),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0  (
    .I(\BU2/U0/TRIMAC_INST_FLOW__n0001 ),
    .CE(\BU2/U0/TRIMAC_INST_FLOW__n0007 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0.GSR.OR ),
    .CLK(txcoreclk),
    .O(emacclienttxstats[31]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG_674 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG_674  (
    .I(\BU2/U0/TRIMAC_INST_FLOW__n0002 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG_675 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG_675  (
    .I(\BU2/U0/TRIMAC_INST_FLOW__n0003 ),
    .RST(\BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [4]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [5]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [4]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [5]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [6]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [7]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [8]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [8]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [9]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [9]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [10]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [10]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [11]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<2>1 .INIT = 16'hEEEB;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_LOAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [1]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [2])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2_676 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2_676  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1_677 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1_677  (
    .I(phyemaccol),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1_678 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1_678  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL_679 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL_679  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0016 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY_680 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY_680  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0015 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY_681 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY_681  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0014 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [7]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2_682 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2_682  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2_683 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2_683  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2_684 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2_684  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1_685 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1_685  (
    .I(\BU2/U0/TRIMAC_INST_INT_EXTENSION ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1_686 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1_686  (
    .I(\BU2/U0/TRIMAC_INST__n0012 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1_687 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1_687  (
    .I(\BU2/U0/TRIMAC_INST__n0011 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [7]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [7]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_GMII_TX_ER_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_GMII_TX_ER_Result1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424_SW0 .INIT = 4'hD;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0424_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START ),
    .O(\BU2/U0/N53281 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068_688 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068_688  (
    .ADR0(\BU2/U0/N65588 ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_N16073 ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [7]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [0]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068 )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068_SW1 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER__n0068_SW1  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7 [3]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL [0]),
    .O(\BU2/U0/N65588 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16_SW0 .INIT = 16'hDC10;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16_SW0  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0183 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0182 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [9]),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_INT_BACK_OFF_TIME [6]),
    .O(\BU2/U0/N65476 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD1 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_N17850 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD1 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_N17850 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_EXTENSION_REG_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_EXTENSION_REG_Result1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_GMII_TX_EN_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Mmux_GMII_TX_EN_Result1  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0059_Result .INIT = 16'hAC5C;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN_Mmux__n0059_Result  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0320 [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE ),
    .ADR3(\BU2/U0/N65768 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRCGEN__n0059 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [6]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL1 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION1 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [3]),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [2]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [5]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [4]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00161 .INIT = 8'h23;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00161  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0016 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0205_Result1 .INIT = 16'h08F8;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_Mmux__n0205_Result1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS ),
    .ADR2(\BU2/U0/N66138 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0205 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<0>1 .INIT = 16'h00F7;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_N17850 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [6]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<1>1 .INIT = 8'h09;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_LOAD ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [3]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [3]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<1>1 .INIT = 8'h09;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<1>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [1]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [1])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<0>1 .INIT = 4'h1;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_261 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_261  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT [4]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_COUNT_inst_lut3_26 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut3 .INIT = 4'h6;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_Eq_stagelut3  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER [8]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_N4293 )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089<15>16  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0224 [15]),
    .ADR1(\BU2/U0/N65478 ),
    .ADR2(\BU2/U0/N65476 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0089 [15])
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Ker178481 .INIT = 8'h08;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_Ker178481  (
    .ADR0(tieemacconfigvec_7[55]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_N17850 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [4]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<0>1 .INIT = 8'h75;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_Mmux__n0001_Result<0>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [0])
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>67_G .INIT = 8'hFB;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX__n0014<7>67_G  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD [39]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT [3]),
    .ADR2(\BU2/U0/CHOICE2875 ),
    .O(\BU2/U0/N66099 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00461 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n00461  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_LOAD ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6  (
    .I(\BU2/U0/TRIMAC_INST__n0009 [6]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0044 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [1]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0046 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00121 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00121  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE ),
    .ADR1(\BU2/U0/CHOICE2257 ),
    .ADR2(\BU2/U0/CHOICE2262 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0012 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7  (
    .I(phyemacrxd_1[7]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [7]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3_689 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3_689  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL_690 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL_690  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0011 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5  (
    .I(phyemacrxd_1[5]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [5]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG_691 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG_691  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_INT_ALIGNMENT_ERR_PULSE ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1_692 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1_692  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0012 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2_693 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2_693  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1_694 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1_694  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2_695 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2_695  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE_696 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE_696  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0020 ),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0054 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE ),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001010 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n001010  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [2]),
    .ADR3(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [3]),
    .O(\BU2/U0/CHOICE3280 )
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001421 .INIT = 16'hFFFE;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE__n001421  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [2]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [4]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX [5]),
    .O(\BU2/U0/CHOICE2045 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2_697 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2_697  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0002 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2_698 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2_698  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR1 .INIT = 8'h80;
  X_LUT3 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR1  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt_699 .INIT = 4'hA;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt_699  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q [5]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CALCULATE_CRC2_CRC1_Q<5>_rt ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004540 .INIT = 16'hF444;
  X_LUT4 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n004540  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_EN_WREN_REG ),
    .ADR1(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR ),
    .ADR2(\BU2/U0/TRIMAC_INST_RXGEN_WR_EN ),
    .ADR3(\BU2/U0/N65759 ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1_700 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1_700  (
    .I(phyemacrxdv),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3_701 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3_701  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0010 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker169021 .INIT = 16'h1000;
  X_LUT4 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_Ker169021  (
    .ADR0(tieemacconfigvec_7[66]),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .ADR3(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_INT_ALIGNMENT_ERR_PULSE )
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04531 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n04531  (
    .ADR0(\BU2/U0/CHOICE2424 ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0315 ),
    .ADR3(\BU2/U0/CHOICE2430 ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0453 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_LPM_COUNTER_14__n0000<0>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_LPM_COUNTER_14__n0000<0>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT [0]),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_N4073 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00201 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n00201  (
    .ADR0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN__n0020 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0  (
    .I(phyemacrxd_1[0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1  (
    .I(phyemacrxd_1[1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3  (
    .I(phyemacrxd_1[3]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [3]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4  (
    .I(phyemacrxd_1[4]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [4]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n045413 .INIT = 16'h0080;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n045413  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0257 ),
    .O(\BU2/U0/CHOICE2655 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2  (
    .I(phyemacrxd_1[2]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [2]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0014 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [1]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [0]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_N4073 ),
    .CE(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2 ),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05261 .INIT = 8'hF2;
  X_LUT3 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n05261  (
    .ADR0(\BU2/U0/TRIMAC_INST_INT_TX_DATA_VALID_OUT ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0526 )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6  (
    .I(phyemacrxd_1[6]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1 [6]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1_702 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1_702  (
    .I(phyemacrxer),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1 ),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<3>1 .INIT = 16'hE000;
  X_LUT4 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151<3>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN ),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN ),
    .ADR2(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1 ),
    .ADR3(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0246 [3]),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1__n0151 [3])
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [1]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [1]),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0002 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [0]),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0016 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY [2]),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [2]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [2]),
    .CE(VCC),
    .SET(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1_703 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1_703 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1_703  (
    .I(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR__n0001 [6]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO__n0045 ),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6.GSR.OR ),
    .SET(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [6])
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT_704 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT_704  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3_705 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3_705  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3 ),
    .CE(VCC),
    .RST(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1_706 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1_706 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1_706  (
    .I(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>lut .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<7>lut  (
    .ADR0(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR [7]),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4378 ),
    .ADR1(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT_707 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT_707  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3_708 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3_708  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3 ),
    .CE(VCC),
    .RST(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1_709 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1_709 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1_709  (
    .I(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1 ),
    .CE(VCC),
    .RST(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<4>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4370 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT_710 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT_710  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3_711 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3_711  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3 ),
    .CE(VCC),
    .RST(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1_712 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1_712 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1_712  (
    .I(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1 ),
    .CE(VCC),
    .RST(GND)
  );
  initial assign \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0 .notifier = 1'bx;
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY [0]),
    .RST(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC [0]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_713 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_713  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3_714 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3_714  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<4>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<4>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [4]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [4]),
    .O(emacphytxd_0[4])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<3>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<3>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [3]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [3]),
    .O(emacphytxd_0[3])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<2>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [2]),
    .O(emacphytxd_0[2])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<1>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<1>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [1]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [1]),
    .O(emacphytxd_0[1])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<0>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<0>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [0]),
    .O(emacphytxd_0[0])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<6>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<6>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [6]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [6]),
    .O(emacphytxd_0[6])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<6>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[6]),
    .ADR2(\BU2/U0/CHOICE2373 ),
    .ADR3(\BU2/U0/N65520 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [6])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<5>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[5]),
    .ADR2(\BU2/U0/CHOICE2349 ),
    .ADR3(\BU2/U0/N65516 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [5])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<4>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[4]),
    .ADR2(\BU2/U0/CHOICE2361 ),
    .ADR3(\BU2/U0/N65512 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [4])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<3>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[3]),
    .ADR2(\BU2/U0/CHOICE2337 ),
    .ADR3(\BU2/U0/N65508 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [3])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<2>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[2]),
    .ADR2(\BU2/U0/CHOICE2313 ),
    .ADR3(\BU2/U0/N65504 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [2])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<1>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[1]),
    .ADR2(\BU2/U0/CHOICE2325 ),
    .ADR3(\BU2/U0/N65500 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [1])
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<0>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[0]),
    .ADR2(\BU2/U0/CHOICE2301 ),
    .ADR3(\BU2/U0/N65496 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [0])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_0 .INIT = 1'b0;
  X_SFF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG_0  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG ),
    .SRST(corehassgmii),
    .SSET(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_INT_ALIGNMENT_ERR_PULSE ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_D_WR_REG [0]),
    .CE(VCC),
    .SET(GND),
    .RST(GSR)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<7>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TXD_Result<7>1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0035 [7]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [7]),
    .O(emacphytxd_0[7])
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR__n0001 [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR [0]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2_715 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2_715  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2.GSR.OR ),
    .CLK(txcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH1  (
    .ADR0(reset),
    .ADR1(tieemacconfigvec_7[60]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH )
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2_716 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2_716  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2_717 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2_717  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2.GSR.OR ),
    .CLK(rxcoreclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR [1]),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2_718 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2_718  (
    .I(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1 ),
    .SET(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2 ),
    .CE(VCC),
    .RST(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<2>1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_FLOW_TX_Mmux_DATA_OUT_Result<2>1  (
    .ADR0(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1 ),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL [2]),
    .ADR2(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT [2]),
    .O(\BU2/U0/TRIMAC_INST_INT_TX_DATA_OUT [2])
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_N4374 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN__n0013 [5]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5.GSR.OR ),
    .CLK(txgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY [5]),
    .CE(VCC),
    .SET(GND)
  );
  X_MUX2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>cy  (
    .IB(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<5>_cyo ),
    .SEL(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_N4374 ),
    .IA(\BU2/U0/address_valid_early ),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_LPM_COUNTER_2__n0004<6>_cyo )
  );
  defparam \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1 .INIT = 1'b0;
  X_FF \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1  (
    .I(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3 [1]),
    .RST(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4 [1]),
    .CE(VCC),
    .SET(GND)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TX_EN_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TX_EN_Result1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0037 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY ),
    .O(emacphytxen)
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_GMII_TX_ER_Result1 .INIT = 8'hD8;
  X_LUT3 \BU2/U0/TRIMAC_INST_Mmux_GMII_TX_ER_Result1  (
    .ADR0(corehassgmii),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN__n0038 [0]),
    .ADR2(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY ),
    .O(emacphytxer)
  );
  defparam \BU2/U0/TRIMAC_INST_FLOW_RX__n00401 .INIT = 16'hFBFA;
  X_LUT4 \BU2/U0/TRIMAC_INST_FLOW_RX__n00401  (
    .ADR0(NlwRenamedSig_OI_emacclientrxstats[0]),
    .ADR1(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT [0]),
    .ADR2(NlwRenamedSig_OI_emacclientrxstats[1]),
    .ADR3(\BU2/U0/TRIMAC_INST_FLOW_RX_N18517 ),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX__n0040 )
  );
  defparam \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>39 .INIT = 16'hDDD8;
  X_LUT4 \BU2/U0/TRIMAC_INST_Mmux_INT_GMII_RXD_Result<7>39  (
    .ADR0(corehassgmii),
    .ADR1(phyemacrxd_1[7]),
    .ADR2(\BU2/U0/CHOICE2289 ),
    .ADR3(\BU2/U0/N65492 ),
    .O(\BU2/U0/TRIMAC_INST_INT_GMII_RXD [7])
  );
  defparam \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_Mmux_WR_OCCUPANCY_Result<1>50  (
    .ADR0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC [0]),
    .ADR1(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR [0]),
    .O(\BU2/U0/CHOICE1724 )
  );
  defparam \BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH1 .INIT = 4'hE;
  X_LUT2 \BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH1  (
    .ADR0(reset),
    .ADR1(tieemacconfigvec_7[53]),
    .O(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH )
  );
  defparam \BU2/U0/TRIMAC_INST__n00031 .INIT = 4'h2;
  X_LUT2 \BU2/U0/TRIMAC_INST__n00031  (
    .ADR0(tieemacconfigvec_7[65]),
    .ADR1(tieemacconfigvec_7[66]),
    .O(speedis100)
  );
  defparam \BU2/U0/TRIMAC_INST_SPEED_IS_10_1001 .INIT = 4'h5;
  X_LUT2 \BU2/U0/TRIMAC_INST_SPEED_IS_10_1001  (
    .ADR0(tieemacconfigvec_7[66]),
    .O(NlwRenamedSig_OI_speedis10100),
    .ADR1(GND)
  );
  X_ONE \BU2/U0/XST_VCC  (
    .O(\BU2/U0/address_valid_early )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2 .INIT = 1'b1;
  X_FF \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2  (
    .I(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR__n0001 [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE ),
    .SET(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2.GSR.OR ),
    .CLK(rxgmiimiiclk),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR [2]),
    .RST(GND)
  );
  X_ZERO \BU2/U0/XST_GND  (
    .O(\NlwRenamedSig_OI_BU2/emacphymclkout )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [7]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN__n0049 ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD7/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [6]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [6]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD6/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [5]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [5]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD5/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [4]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [4]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD4/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [3]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [3]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD3/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [2]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [2]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD2/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [1]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [1]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD1/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1 [0]),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG5 [0]),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RXD0/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG5 ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_DV/SRL16E_Q15_UNCONNECTED )
  );
  X_ONE \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/VCC  (
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/CE )
  );
  defparam \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/SRL16E .INIT = 16'h0000;
  X_SRLC16E \BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/SRL16E  (
    .D(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1 ),
    .CE(\BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/CE ),
    .CLK(rxcoreclk),
    .A3(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A2(\NlwRenamedSig_OI_BU2/emacphymclkout ),
    .A1(\BU2/U0/address_valid_early ),
    .A0(\BU2/U0/address_valid_early ),
    .Q(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG5 ),
    .Q15(\NLW_BU2/U0/TRIMAC_INST_RXGEN_DELAY_RX_ERR/SRL16E_Q15_UNCONNECTED )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7.GSR.OR_719  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6.GSR.OR_720  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5.GSR.OR_721  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4.GSR.OR_722  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3.GSR.OR_723  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2.GSR.OR_724  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1.GSR.OR_725  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1.GSR.OR_726  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1.GSR.OR_727  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1.GSR.OR_728  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1.GSR.OR_729  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1.GSR.OR_730  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG.GSR.OR_731  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_MIFG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE.GSR.OR_732  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1.GSR.OR_733  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0.GSR.OR_734  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0.GSR.OR_735  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE.GSR.OR_736  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR.GSR.OR_737  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MAX_LENGTH_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR.GSR.OR_738  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FRAME_LEN_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN.GSR.OR_739  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_EXCEEDED_MIN_LEN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH.GSR.OR_740  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_MIN_LENGTH_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME.GSR.OR_741  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_INHIBIT_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR.GSR.OR_742  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT.GSR.OR_743  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_ALIGNMENT_ERROR_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR.GSR.OR_744  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_OUT_OF_BOUNDS_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR.GSR.OR_745  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_CRC_ENGINE_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME.GSR.OR_746  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_BAD_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME.GSR.OR_747  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_GOOD_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID.GSR.OR_748  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_STATISTICS_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR.GSR.OR_749  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_FCS_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44.GSR.OR_750  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_44.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43.GSR.OR_751  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_43.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12.GSR.OR_752  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11.GSR.OR_753  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10.GSR.OR_754  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9.GSR.OR_755  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8.GSR.OR_756  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7.GSR.OR_757  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6.GSR.OR_758  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5.GSR.OR_759  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4.GSR.OR_760  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3.GSR.OR_761  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2.GSR.OR_762  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1.GSR.OR_763  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0.GSR.OR_764  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41.GSR.OR_765  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_41.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39.GSR.OR_766  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_39.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID.GSR.OR_767  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS.GSR.OR_768  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_NO_FCS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS.GSR.OR_769  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_WITH_FCS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME.GSR.OR_770  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_PADDED_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE.GSR.OR_771  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ONE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO.GSR.OR_772  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_ZERO.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256.GSR.OR_773  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LESS_THAN_256.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH.GSR.OR_774  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0.GSR.OR_775  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1.GSR.OR_776  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2.GSR.OR_777  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3.GSR.OR_778  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4.GSR.OR_779  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5.GSR.OR_780  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6.GSR.OR_781  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7.GSR.OR_782  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8.GSR.OR_783  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9.GSR.OR_784  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10.GSR.OR_785  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_DATA_COUNTER_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0.GSR.OR_786  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1.GSR.OR_787  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2.GSR.OR_788  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3.GSR.OR_789  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4.GSR.OR_790  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5.GSR.OR_791  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6.GSR.OR_792  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7.GSR.OR_793  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8.GSR.OR_794  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9.GSR.OR_795  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10.GSR.OR_796  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_LENGTH_TYPE_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE.GSR.OR_797  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CRC_COMPUTE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET.GSR.OR_798  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_TYPE_PACKET.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5.GSR.OR_799  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4.GSR.OR_800  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3.GSR.OR_801  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2.GSR.OR_802  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1.GSR.OR_803  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0.GSR.OR_804  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_PAUSE_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5.GSR.OR_805  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4.GSR.OR_806  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3.GSR.OR_807  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2.GSR.OR_808  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1.GSR.OR_809  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0.GSR.OR_810  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADDRESS_MATCH_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH.GSR.OR_811  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE.GSR.OR_812  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT.GSR.OR_813  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME.GSR.OR_814  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_ADD_CONTROL_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42.GSR.OR_815  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_42.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38.GSR.OR_816  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_38.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40.GSR.OR_817  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_40.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30.GSR.OR_818  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_30.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31.GSR.OR_819  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_31.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32.GSR.OR_820  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_32.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33.GSR.OR_821  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_33.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34.GSR.OR_822  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_34.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35.GSR.OR_823  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_35.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36.GSR.OR_824  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_36.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37.GSR.OR_825  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_FRAME_COUNTER_37.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13.GSR.OR_826  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_STATISTICS_LENGTH_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG.GSR.OR_827  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_RX_DV_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH.GSR.OR_828  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME.GSR.OR_829  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_MULTICAST_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME.GSR.OR_830  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5.GSR.OR_831  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4.GSR.OR_832  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3.GSR.OR_833  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2.GSR.OR_834  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1.GSR.OR_835  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0.GSR.OR_836  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_BROADCAST_MATCH_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH.GSR.OR_837  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME.GSR.OR_838  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_VLAN_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT.GSR.OR_839  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME.GSR.OR_840  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_DECODER_CONTROL_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME.GSR.OR_841  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_FRAME.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE.GSR.OR_842  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_PREAMBLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD.GSR.OR_843  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DAT_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA.GSR.OR_844  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_END_DATA.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD.GSR.OR_845  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_DEST_ADDRESS_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD.GSR.OR_846  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_SRC_ADDRESS_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD.GSR.OR_847  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_CRC_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD.GSR.OR_848  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_EXT_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5.GSR.OR_849  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4.GSR.OR_850  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3.GSR.OR_851  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2.GSR.OR_852  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1.GSR.OR_853  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0.GSR.OR_854  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_FIELD_CONTROL_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG.GSR.OR_855  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_DV_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC.GSR.OR_856  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_RATE_GEN_SYNC.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42.GSR.OR_857  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_42.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41.GSR.OR_858  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_41.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40.GSR.OR_859  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_40.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39.GSR.OR_860  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_39.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38.GSR.OR_861  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_38.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37.GSR.OR_862  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_37.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36.GSR.OR_863  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_36.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35.GSR.OR_864  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_35.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34.GSR.OR_865  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_34.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33.GSR.OR_866  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_33.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32.GSR.OR_867  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_32.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31.GSR.OR_868  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_31.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30.GSR.OR_869  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_30.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29.GSR.OR_870  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_29.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28.GSR.OR_871  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_28.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27.GSR.OR_872  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_27.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26.GSR.OR_873  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_26.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25.GSR.OR_874  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_25.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24.GSR.OR_875  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_24.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23.GSR.OR_876  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_23.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22.GSR.OR_877  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_22.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21.GSR.OR_878  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_21.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20.GSR.OR_879  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_20.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19.GSR.OR_880  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_19.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18.GSR.OR_881  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17.GSR.OR_882  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16.GSR.OR_883  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15.GSR.OR_884  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14.GSR.OR_885  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13.GSR.OR_886  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12.GSR.OR_887  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11.GSR.OR_888  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10.GSR.OR_889  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9.GSR.OR_890  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8.GSR.OR_891  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7.GSR.OR_892  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6.GSR.OR_893  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5.GSR.OR_894  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4.GSR.OR_895  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3.GSR.OR_896  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2.GSR.OR_897  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1.GSR.OR_898  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0.GSR.OR_899  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6.GSR.OR_900  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5.GSR.OR_901  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4.GSR.OR_902  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3.GSR.OR_903  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2.GSR.OR_904  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1.GSR.OR_905  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0.GSR.OR_906  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6.GSR.OR_907  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5.GSR.OR_908  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4.GSR.OR_909  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3.GSR.OR_910  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2.GSR.OR_911  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1.GSR.OR_912  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0.GSR.OR_913  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6.GSR.OR_914  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5.GSR.OR_915  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4.GSR.OR_916  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3.GSR.OR_917  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2.GSR.OR_918  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1.GSR.OR_919  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0.GSR.OR_920  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6.GSR.OR_921  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5.GSR.OR_922  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4.GSR.OR_923  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3.GSR.OR_924  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2.GSR.OR_925  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1.GSR.OR_926  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0.GSR.OR_927  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6.GSR.OR_928  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5.GSR.OR_929  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4.GSR.OR_930  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3.GSR.OR_931  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2.GSR.OR_932  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1.GSR.OR_933  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0.GSR.OR_934  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_6.GSR.OR_935  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_5.GSR.OR_936  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_4.GSR.OR_937  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_3.GSR.OR_938  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_2.GSR.OR_939  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_1.GSR.OR_940  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_0.GSR.OR_941  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD.GSR.OR_942  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_LT_CHECK_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD.GSR.OR_943  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_HALF_DUPLEX_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD.GSR.OR_944  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CRC_MODE_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD.GSR.OR_945  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_VLAN_ENABLE_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD.GSR.OR_946  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_JUMBO_FRAMES_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47.GSR.OR_947  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_47.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG.GSR.OR_948  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_ENABLE_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0.GSR.OR_949  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1.GSR.OR_950  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2.GSR.OR_951  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3.GSR.OR_952  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4.GSR.OR_953  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5.GSR.OR_954  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6.GSR.OR_955  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7.GSR.OR_956  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8.GSR.OR_957  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9.GSR.OR_958  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10.GSR.OR_959  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11.GSR.OR_960  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12.GSR.OR_961  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13.GSR.OR_962  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14.GSR.OR_963  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15.GSR.OR_964  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16.GSR.OR_965  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17.GSR.OR_966  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18.GSR.OR_967  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19.GSR.OR_968  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_19.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20.GSR.OR_969  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_20.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21.GSR.OR_970  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_21.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22.GSR.OR_971  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_22.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23.GSR.OR_972  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_23.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24.GSR.OR_973  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VECTOR_24.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG.GSR.OR_974  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_ALIGNMENT_ERROR_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID.GSR.OR_975  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_STATISTICS_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT.GSR.OR_976  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG5_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT.GSR.OR_977  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG4_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT.GSR.OR_978  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG3_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT.GSR.OR_979  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG2_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT.GSR.OR_980  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_CE_REG1_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT.GSR.OR_981  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG5_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT.GSR.OR_982  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG4_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT.GSR.OR_983  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG3_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT.GSR.OR_984  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG2_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT.GSR.OR_985  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_REG1_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR.GSR.OR_986  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_FRAME_CHECKER_SLOT_LENGTH_ERROR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD.GSR.OR_987  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_SM_LEN_FIELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7.GSR.OR_988  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG8_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_7.GSR.OR_989  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG.GSR.OR_990  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SFD_FLAG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG.GSR.OR_991  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_EXTENSION_FLAG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD.GSR.OR_992  (
    .I0(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_SPEED_IS_10_100_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7.GSR.OR_993  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_WR_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43.GSR.OR_994  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_43.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR.GSR.OR_995  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_WR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR.GSR.OR_996  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_WR.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1.GSR.OR_997  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2.GSR.OR_998  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44.GSR.OR_999  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_44.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46.GSR.OR_1000  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_46.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45.GSR.OR_1001  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_PAUSE_ADD_HELD_45.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6.GSR.OR_1002  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7.GSR.OR_1003  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_DV_REG7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1.GSR.OR_1004  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6.GSR.OR_1005  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7.GSR.OR_1006  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_ERR_REG7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7.GSR.OR_1007  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG1_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7.GSR.OR_1008  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG6_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7.GSR.OR_1009  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RXD_REG7_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0.GSR.OR_1010  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1.GSR.OR_1011  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID.GSR.OR_1012  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_DATA_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1.GSR.OR_1013  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0.GSR.OR_1014  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1.GSR.OR_1015  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2.GSR.OR_1016  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0.GSR.OR_1017  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6.GSR.OR_1018  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_6__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7.GSR.OR_1019  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_7__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0.GSR.OR_1020  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_0__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2.GSR.OR_1021  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2.GSR.OR_1022  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_2__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5.GSR.OR_1023  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_5__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4.GSR.OR_1024  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_4__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3.GSR.OR_1025  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_3__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1.GSR.OR_1026  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2.GSR.OR_1027  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1.GSR.OR_1028  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0.GSR.OR_1029  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDRGRAY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2.GSR.OR_1030  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2.GSR.OR_1031  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1.GSR.OR_1032  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0.GSR.OR_1033  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDRGRAY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0.GSR.OR_1034  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1.GSR.OR_1035  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RAG_WRITESYNC_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2.GSR.OR_1036  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_RD_ADDR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1.GSR.OR_1037  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_0_1__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_IFG_CNTR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1.GSR.OR_1038  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WAG_READSYNC_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG.GSR.OR_1039  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_MIFG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE.GSR.OR_1040  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1.GSR.OR_1041  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0.GSR.OR_1042  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_NEXT_WR_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0.GSR.OR_1043  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_WR_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE.GSR.OR_1044  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5.GSR.OR_1045  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1.GSR.OR_1046  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2.GSR.OR_1047  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1.GSR.OR_1048  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3.GSR.OR_1049  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2.GSR.OR_1050  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0.GSR.OR_1051  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_IFG_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3.GSR.OR_1052  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4.GSR.OR_1053  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5.GSR.OR_1054  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6.GSR.OR_1055  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1.GSR.OR_1056  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15.GSR.OR_1057  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14.GSR.OR_1058  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13.GSR.OR_1059  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12.GSR.OR_1060  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11.GSR.OR_1061  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10.GSR.OR_1062  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9.GSR.OR_1063  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8.GSR.OR_1064  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7.GSR.OR_1065  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6.GSR.OR_1066  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5.GSR.OR_1067  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4.GSR.OR_1068  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3.GSR.OR_1069  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2.GSR.OR_1070  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1.GSR.OR_1071  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0.GSR.OR_1072  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17.GSR.OR_1073  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18.GSR.OR_1074  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4.GSR.OR_1075  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1.GSR.OR_1076  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5.GSR.OR_1077  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0.GSR.OR_1078  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1.GSR.OR_1079  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2.GSR.OR_1080  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3.GSR.OR_1081  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2.GSR.OR_1082  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_MAX_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4.GSR.OR_1083  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6.GSR.OR_1084  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7.GSR.OR_1085  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8.GSR.OR_1086  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11.GSR.OR_1087  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10.GSR.OR_1088  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3.GSR.OR_1089  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8.GSR.OR_1090  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8.GSR.OR_1091  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7.GSR.OR_1092  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0.GSR.OR_1093  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7.GSR.OR_1094  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1.GSR.OR_1095  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2.GSR.OR_1096  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6.GSR.OR_1097  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0.GSR.OR_1098  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1.GSR.OR_1099  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0.GSR.OR_1100  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1.GSR.OR_1101  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0.GSR.OR_1102  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7.GSR.OR_1103  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12.GSR.OR_1104  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10.GSR.OR_1105  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4.GSR.OR_1106  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3.GSR.OR_1107  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0001 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1.GSR.OR_1108  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0.GSR.OR_1109  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13.GSR.OR_1110  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14.GSR.OR_1111  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_3__n0001 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER_COUNT_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6.GSR.OR_1112  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10.GSR.OR_1113  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8.GSR.OR_1114  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5.GSR.OR_1115  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9.GSR.OR_1116  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10.GSR.OR_1117  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11.GSR.OR_1118  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3.GSR.OR_1119  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12.GSR.OR_1120  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13.GSR.OR_1121  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14.GSR.OR_1122  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15.GSR.OR_1123  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16.GSR.OR_1124  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2.GSR.OR_1125  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17.GSR.OR_1126  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18.GSR.OR_1127  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19.GSR.OR_1128  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_19.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID.GSR.OR_1129  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20.GSR.OR_1130  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_20.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE.GSR.OR_1131  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DEFER_COUNT_DONE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12.GSR.OR_1132  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED.GSR.OR_1133  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2.GSR.OR_1134  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DEFERRED2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET.GSR.OR_1135  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_QUIET.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS.GSR.OR_1136  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_CRS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID.GSR.OR_1137  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_DATA_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION.GSR.OR_1138  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_LATE_COLLISION.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS.GSR.OR_1139  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_EXCESSIVE_COLLISIONS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3.GSR.OR_1140  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT.GSR.OR_1141  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_MAX_PKT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH.GSR.OR_1142  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_SCSH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21.GSR.OR_1143  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_21.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22.GSR.OR_1144  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_22.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14.GSR.OR_1145  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN.GSR.OR_1146  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_VLAN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL.GSR.OR_1147  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_CONTROL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15.GSR.OR_1148  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH.GSR.OR_1149  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE5_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH.GSR.OR_1150  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_MULTI_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH.GSR.OR_1151  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE4_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH.GSR.OR_1152  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE3_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH.GSR.OR_1153  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE2_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH.GSR.OR_1154  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE1_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH.GSR.OR_1155  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DST_ADDR_BYTE0_MATCH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS.GSR.OR_1156  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_SUCCESS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2.GSR.OR_1157  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN.GSR.OR_1158  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_UNDERRUN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID.GSR.OR_1159  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_STATUS_VALID.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL.GSR.OR_1160  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_COL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT.GSR.OR_1161  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_RETRANSMIT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START.GSR.OR_1162  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_START.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX.GSR.OR_1163  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CR178124_FIX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0.GSR.OR_1164  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD_PIPE_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0.GSR.OR_1165  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1.GSR.OR_1166  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT_PIPE_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1.GSR.OR_1167  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2.GSR.OR_1168  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3.GSR.OR_1169  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4.GSR.OR_1170  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5.GSR.OR_1171  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6.GSR.OR_1172  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7.GSR.OR_1173  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8.GSR.OR_1174  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9.GSR.OR_1175  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10.GSR.OR_1176  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11.GSR.OR_1177  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12.GSR.OR_1178  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13.GSR.OR_1179  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE_PIPE_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7.GSR.OR_1180  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7.GSR.OR_1181  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7.GSR.OR_1182  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7.GSR.OR_1183  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7.GSR.OR_1184  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE.GSR.OR_1185  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COMPUTE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION.GSR.OR_1186  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_EXTENSION.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC.GSR.OR_1187  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD.GSR.OR_1188  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PAD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT.GSR.OR_1189  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TRANSMIT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE.GSR.OR_1190  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE.GSR.OR_1191  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PREAMBLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER.GSR.OR_1192  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DEFER.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY.GSR.OR_1193  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_PRE_DELAY.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN.GSR.OR_1194  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF_SEEN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23.GSR.OR_1195  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_23.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED.GSR.OR_1196  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MAX_PKT_LEN_REACHED.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED.GSR.OR_1197  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIN_PKT_LEN_REACHED.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED.GSR.OR_1198  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SLOT_TIME_REACHED.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16.GSR.OR_1199  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BACK_OFF_COUNT_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0.GSR.OR_1200  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1.GSR.OR_1201  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3.GSR.OR_1202  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE.GSR.OR_1203  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_PREAMBLE_DONE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2.GSR.OR_1204  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL.GSR.OR_1205  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_FAIL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL.GSR.OR_1206  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_EARLY_COL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL.GSR.OR_1207  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_COL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT.GSR.OR_1208  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_WFBOT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED.GSR.OR_1209  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COL_SAVED.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM.GSR.OR_1210  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_JAM.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH.GSR.OR_1211  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_MAX_LENGTH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER.GSR.OR_1212  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BURST_OVER.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE.GSR.OR_1213  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CLIENT_FRAME_DONE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG.GSR.OR_1214  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_MIFG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG.GSR.OR_1215  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETIFG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST.GSR.OR_1216  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETST.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK.GSR.OR_1217  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX_OK.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH.GSR.OR_1218  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_ETSCSH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD.GSR.OR_1219  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_BAD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD.GSR.OR_1220  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FRAME_GOOD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH.GSR.OR_1221  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_SCSH.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS.GSR.OR_1222  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_FCS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF.GSR.OR_1223  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_COF.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL.GSR.OR_1224  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CFL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA.GSR.OR_1225  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_DA.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX.GSR.OR_1226  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_TX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE.GSR.OR_1227  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS.GSR.OR_1228  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CDS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL.GSR.OR_1229  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IDL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7.GSR.OR_1230  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7.GSR.OR_1231  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100.GSR.OR_1232  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100__n0000 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_SPEED_IS_10_100.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7.GSR.OR_1233  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7.GSR.OR_1234  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN.GSR.OR_1235  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX.GSR.OR_1236  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_HALF_DUPLEX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN.GSR.OR_1237  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_VLAN_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN.GSR.OR_1238  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_JUMBO_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE.GSR.OR_1239  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_CRC_MODE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1.GSR.OR_1240  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN.GSR.OR_1241  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_EN_IN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4.GSR.OR_1242  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6.GSR.OR_1243  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5.GSR.OR_1244  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4.GSR.OR_1245  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0.GSR.OR_1246  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1.GSR.OR_1247  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2.GSR.OR_1248  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2.GSR.OR_1249  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9.GSR.OR_1250  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3.GSR.OR_1251  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION.GSR.OR_1252  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STOP_EXTENSION.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9.GSR.OR_1253  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6.GSR.OR_1254  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_4_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25.GSR.OR_1255  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_25.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3.GSR.OR_1256  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4.GSR.OR_1257  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2.GSR.OR_1258  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6.GSR.OR_1259  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4.GSR.OR_1260  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3.GSR.OR_1261  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5.GSR.OR_1262  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3.GSR.OR_1263  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14.GSR.OR_1264  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4.GSR.OR_1265  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1.GSR.OR_1266  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5.GSR.OR_1267  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13.GSR.OR_1268  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5.GSR.OR_1269  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2.GSR.OR_1270  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3.GSR.OR_1271  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6.GSR.OR_1272  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5.GSR.OR_1273  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0.GSR.OR_1274  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2.GSR.OR_1275  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_TX_ATTEMPTS_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2.GSR.OR_1276  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3.GSR.OR_1277  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6.GSR.OR_1278  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6.GSR.OR_1279  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0.GSR.OR_1280  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_CRC_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0.GSR.OR_1281  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2.GSR.OR_1282  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1.GSR.OR_1283  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12.GSR.OR_1284  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13.GSR.OR_1285  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0.GSR.OR_1286  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2.GSR.OR_1287  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11.GSR.OR_1288  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1.GSR.OR_1289  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0.GSR.OR_1290  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_PRE_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4.GSR.OR_1291  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6.GSR.OR_1292  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11.GSR.OR_1293  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2.GSR.OR_1294  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6.GSR.OR_1295  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0.GSR.OR_1296  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1.GSR.OR_1297  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0.GSR.OR_1298  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6.GSR.OR_1299  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5.GSR.OR_1300  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_2_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9.GSR.OR_1301  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2.GSR.OR_1302  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0.GSR.OR_1303  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1.GSR.OR_1304  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2.GSR.OR_1305  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2.GSR.OR_1306  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3.GSR.OR_1307  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3.GSR.OR_1308  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4.GSR.OR_1309  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5.GSR.OR_1310  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4.GSR.OR_1311  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_IFG_DELAY_HELD_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1.GSR.OR_1312  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4.GSR.OR_1313  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5.GSR.OR_1314  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3.GSR.OR_1315  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6.GSR.OR_1316  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7.GSR.OR_1317  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8.GSR.OR_1318  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9.GSR.OR_1319  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3.GSR.OR_1320  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10.GSR.OR_1321  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2.GSR.OR_1322  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_CONST_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5.GSR.OR_1323  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LEN_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12.GSR.OR_1324  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4.GSR.OR_1325  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_1_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13.GSR.OR_1326  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_2_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0.GSR.OR_1327  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1.GSR.OR_1328  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2.GSR.OR_1329  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3.GSR.OR_1330  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0.GSR.OR_1331  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_3_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4.GSR.OR_1332  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5.GSR.OR_1333  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_LATE_COUNT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5.GSR.OR_1334  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1.GSR.OR_1335  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6.GSR.OR_1336  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7.GSR.OR_1337  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8.GSR.OR_1338  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9.GSR.OR_1339  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_8 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10.GSR.OR_1340  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11.GSR.OR_1341  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12.GSR.OR_1342  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13.GSR.OR_1343  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_1_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8.GSR.OR_1344  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2.GSR.OR_1345  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0.GSR.OR_1346  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1.GSR.OR_1347  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_9 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_BYTE_COUNT_0_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4.GSR.OR_1348  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3.GSR.OR_1349  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_DATA_REG_0_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1.GSR.OR_1350  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26.GSR.OR_1351  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_26.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2.GSR.OR_1352  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4.GSR.OR_1353  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5.GSR.OR_1354  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DEL_MASKED_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27.GSR.OR_1355  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_27.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN.GSR.OR_1356  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_REG_TX_ER_IN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28.GSR.OR_1357  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_STATUS_VECTOR_28.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5.GSR.OR_1358  (
    .I0(\BU2/U0/TRIMAC_INST_TXGEN_RESETb1_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM1_INT_IFG_DELAY_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1.GSR.OR_1359  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0.GSR.OR_1360  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3.GSR.OR_1361  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4.GSR.OR_1362  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5.GSR.OR_1363  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6.GSR.OR_1364  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7.GSR.OR_1365  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8.GSR.OR_1366  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2.GSR.OR_1367  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9.GSR.OR_1368  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_BOC_Q_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0.GSR.OR_1369  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2.GSR.OR_1370  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1.GSR.OR_1371  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3.GSR.OR_1372  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM3_TX_STATE_FFd3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT.GSR.OR_1373  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG2_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT.GSR.OR_1374  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG1_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4.GSR.OR_1375  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_1 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_SM2_TX_STATE_FFd4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN.GSR.OR_1376  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRC100_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT.GSR.OR_1377  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG1_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT.GSR.OR_1378  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG2_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT.GSR.OR_1379  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG3_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT.GSR.OR_1380  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG4_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT.GSR.OR_1381  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CE_REG5_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT.GSR.OR_1382  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG3_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT.GSR.OR_1383  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG4_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1.GSR.OR_1384  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT.GSR.OR_1385  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_REG5_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG.GSR.OR_1386  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV10_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0.GSR.OR_1387  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_TX_FIFO_RD_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN.GSR.OR_1388  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CRC1000_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_CRS.GSR.OR_1389  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRS.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE.GSR.OR_1390  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_CRC_MODE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX.GSR.OR_1391  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_HALF_DUPLEX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100.GSR.OR_1392  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_SPEED_IS_10_100.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE.GSR.OR_1393  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_JUMBO_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE.GSR.OR_1394  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE.GSR.OR_1395  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_VLAN_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN.GSR.OR_1396  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_INT_IFG_DEL_EN.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES.GSR.OR_1397  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_2 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_NUMBER_OF_BYTES.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG.GSR.OR_1398  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_TXGEN_CLK_DIV100_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6.GSR.OR_1399  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5.GSR.OR_1400  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4.GSR.OR_1401  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3.GSR.OR_1402  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2.GSR.OR_1403  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1.GSR.OR_1404  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0.GSR.OR_1405  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14.GSR.OR_1406  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13.GSR.OR_1407  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12.GSR.OR_1408  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11.GSR.OR_1409  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10.GSR.OR_1410  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9.GSR.OR_1411  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8.GSR.OR_1412  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7.GSR.OR_1413  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6.GSR.OR_1414  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5.GSR.OR_1415  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4.GSR.OR_1416  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3.GSR.OR_1417  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2.GSR.OR_1418  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1.GSR.OR_1419  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0.GSR.OR_1420  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2.GSR.OR_1421  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1.GSR.OR_1422  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0.GSR.OR_1423  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3.GSR.OR_1424  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4.GSR.OR_1425  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25.GSR.OR_1426  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_25.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28.GSR.OR_1427  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_28.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27.GSR.OR_1428  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_27.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30.GSR.OR_1429  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_30.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29.GSR.OR_1430  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_29.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15.GSR.OR_1431  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14.GSR.OR_1432  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23.GSR.OR_1433  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_23.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22.GSR.OR_1434  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_22.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21.GSR.OR_1435  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_21.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31.GSR.OR_1436  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_31.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6.GSR.OR_1437  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24.GSR.OR_1438  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_24.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46.GSR.OR_1439  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_46.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2.GSR.OR_1440  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26.GSR.OR_1441  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_26.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG.GSR.OR_1442  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3.GSR.OR_1443  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_STATE_COUNT_FFd3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT.GSR.OR_1444  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47.GSR.OR_1445  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_47.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11.GSR.OR_1446  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD.GSR.OR_1447  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_END_OF_TX_HELD.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5.GSR.OR_1448  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4.GSR.OR_1449  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1.GSR.OR_1450  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0.GSR.OR_1451  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7.GSR.OR_1452  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2.GSR.OR_1453  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8.GSR.OR_1454  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3.GSR.OR_1455  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9.GSR.OR_1456  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10.GSR.OR_1457  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41.GSR.OR_1458  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_41.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40.GSR.OR_1459  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_40.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39.GSR.OR_1460  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_39.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42.GSR.OR_1461  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_42.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12.GSR.OR_1462  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34.GSR.OR_1463  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_34.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17.GSR.OR_1464  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36.GSR.OR_1465  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_36.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16.GSR.OR_1466  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20.GSR.OR_1467  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_20.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35.GSR.OR_1468  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_35.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43.GSR.OR_1469  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_43.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18.GSR.OR_1470  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44.GSR.OR_1471  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_44.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37.GSR.OR_1472  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_37.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13.GSR.OR_1473  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38.GSR.OR_1474  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_38.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19.GSR.OR_1475  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_19.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45.GSR.OR_1476  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_45.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32.GSR.OR_1477  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_32.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15.GSR.OR_1478  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_VALUE_HELD_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT.GSR.OR_1479  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_REQ_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT.GSR.OR_1480  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ACK_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1.GSR.OR_1481  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7.GSR.OR_1482  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_7 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_CONTROL_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33.GSR.OR_1483  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_4 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_SOURCE_HELD_33.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL.GSR.OR_1484  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_MUX_CONTROL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL.GSR.OR_1485  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_CONTROL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG.GSR.OR_1486  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_AVAIL_IN_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7.GSR.OR_1487  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3.GSR.OR_1488  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4.GSR.OR_1489  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5.GSR.OR_1490  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6.GSR.OR_1491  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7.GSR.OR_1492  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8.GSR.OR_1493  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9.GSR.OR_1494  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10.GSR.OR_1495  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11.GSR.OR_1496  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12.GSR.OR_1497  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13.GSR.OR_1498  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14.GSR.OR_1499  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15.GSR.OR_1500  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT.GSR.OR_1501  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_OPCODE_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT.GSR.OR_1502  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_REQ_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2.GSR.OR_1503  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4.GSR.OR_1504  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1.GSR.OR_1505  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3.GSR.OR_1506  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0.GSR.OR_1507  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2.GSR.OR_1508  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1.GSR.OR_1509  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0.GSR.OR_1510  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_VALUE_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6.GSR.OR_1511  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17.GSR.OR_1512  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_17.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21.GSR.OR_1513  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_21.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20.GSR.OR_1514  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_20.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3.GSR.OR_1515  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2.GSR.OR_1516  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1.GSR.OR_1517  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0.GSR.OR_1518  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18.GSR.OR_1519  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_18.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5.GSR.OR_1520  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13.GSR.OR_1521  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12.GSR.OR_1522  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG.GSR.OR_1523  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9.GSR.OR_1524  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10.GSR.OR_1525  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14.GSR.OR_1526  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15.GSR.OR_1527  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11.GSR.OR_1528  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16.GSR.OR_1529  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_16.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19.GSR.OR_1530  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_19.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET.GSR.OR_1531  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG.GSR.OR_1532  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_COUNT_SET_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX.GSR.OR_1533  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_GOOD_FRAME_IN_TX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8.GSR.OR_1534  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT.GSR.OR_1535  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_STATUS_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4.GSR.OR_1536  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_5 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_QUANTA_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13.GSR.OR_1537  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_13.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12.GSR.OR_1538  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_12.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11.GSR.OR_1539  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10.GSR.OR_1540  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9.GSR.OR_1541  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8.GSR.OR_1542  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7.GSR.OR_1543  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6.GSR.OR_1544  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5.GSR.OR_1545  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4.GSR.OR_1546  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3.GSR.OR_1547  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2.GSR.OR_1548  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1.GSR.OR_1549  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0.GSR.OR_1550  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX.GSR.OR_1551  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_REQ_TO_TX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15.GSR.OR_1552  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_15.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX.GSR.OR_1553  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_TO_TX.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3.GSR.OR_1554  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2.GSR.OR_1555  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1.GSR.OR_1556  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_GOOD_FRAME_IN1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4.GSR.OR_1557  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3.GSR.OR_1558  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2.GSR.OR_1559  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1.GSR.OR_1560  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0.GSR.OR_1561  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6.GSR.OR_1562  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5.GSR.OR_1563  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4.GSR.OR_1564  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3.GSR.OR_1565  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2.GSR.OR_1566  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1.GSR.OR_1567  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0.GSR.OR_1568  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT.GSR.OR_1569  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_BAD_FRAME_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT.GSR.OR_1570  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_GOOD_FRAME_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT.GSR.OR_1571  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_VALID_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7.GSR.OR_1572  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7.GSR.OR_1573  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_PAUSE_PAUSE_COUNT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14.GSR.OR_1574  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_PAUSE_PAUSE_VALUE_TO_TX_14.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7.GSR.OR_1575  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_DATA_INT_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5.GSR.OR_1576  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT.GSR.OR_1577  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_UNDERRUN_INT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6.GSR.OR_1578  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_DATA_INT_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT.GSR.OR_1579  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_3 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_RETRANSMIT_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT.GSR.OR_1580  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_COLLISION_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0.GSR.OR_1581  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_PAUSE_VECTOR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG.GSR.OR_1582  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_RX_ENABLE_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG.GSR.OR_1583  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT_6 ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_FLOW_TX_ENABLE_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3.GSR.OR_1584  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2.GSR.OR_1585  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3.GSR.OR_1586  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4.GSR.OR_1587  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5.GSR.OR_1588  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3.GSR.OR_1589  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3.GSR.OR_1590  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2.GSR.OR_1591  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3.GSR.OR_1592  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4.GSR.OR_1593  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5.GSR.OR_1594  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6.GSR.OR_1595  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7.GSR.OR_1596  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8.GSR.OR_1597  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_8.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9.GSR.OR_1598  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_9.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10.GSR.OR_1599  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_10.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11.GSR.OR_1600  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_11.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2.GSR.OR_1601  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2.GSR.OR_1602  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1.GSR.OR_1603  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_COL_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3.GSR.OR_1604  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1.GSR.OR_1605  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL.GSR.OR_1606  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_MUXSEL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY.GSR.OR_1607  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_ER_TO_PHY.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY.GSR.OR_1608  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TX_EN_TO_PHY.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7.GSR.OR_1609  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2.GSR.OR_1610  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2.GSR.OR_1611  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2.GSR.OR_1612  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1.GSR.OR_1613  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_EXTENSION_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1.GSR.OR_1614  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_ER_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1.GSR.OR_1615  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TX_EN_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7.GSR.OR_1616  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7.GSR.OR_1617  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1.GSR.OR_1618  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0.GSR.OR_1619  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_DELAY_SHIFT_REG_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2.GSR.OR_1620  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6.GSR.OR_1621  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5.GSR.OR_1622  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1.GSR.OR_1623  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4.GSR.OR_1624  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0.GSR.OR_1625  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1.GSR.OR_1626  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6.GSR.OR_1627  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3.GSR.OR_1628  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1.GSR.OR_1629  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0.GSR.OR_1630  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0.GSR.OR_1631  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1.GSR.OR_1632  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4.GSR.OR_1633  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0.GSR.OR_1634  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG2_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6.GSR.OR_1635  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_TXD_REG1_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2.GSR.OR_1636  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_PREAMBLE_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0.GSR.OR_1637  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1.GSR.OR_1638  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2.GSR.OR_1639  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_NORMAL_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0.GSR.OR_1640  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1.GSR.OR_1641  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2.GSR.OR_1642  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_JAM_EXTENSION_COUNT_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2.GSR.OR_1643  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3.GSR.OR_1644  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0.GSR.OR_1645  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1.GSR.OR_1646  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2.GSR.OR_1647  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3.GSR.OR_1648  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG3_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0.GSR.OR_1649  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1.GSR.OR_1650  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2.GSR.OR_1651  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3.GSR.OR_1652  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG2_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7.GSR.OR_1653  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_7.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3.GSR.OR_1654  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL.GSR.OR_1655  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_MUXSEL.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5.GSR.OR_1656  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG.GSR.OR_1657  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_ALIGNMENT_ERR_REG.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1.GSR.OR_1658  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2.GSR.OR_1659  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_COMB_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1.GSR.OR_1660  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2.GSR.OR_1661  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_NO_ERROR_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE.GSR.OR_1662  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2.GSR.OR_1663  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2.GSR.OR_1664  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0.GSR.OR_1665  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2.GSR.OR_1666  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1.GSR.OR_1667  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3.GSR.OR_1668  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_DV_REG3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0.GSR.OR_1669  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1.GSR.OR_1670  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3.GSR.OR_1671  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4.GSR.OR_1672  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_4.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2.GSR.OR_1673  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1.GSR.OR_1674  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RD_ADDRGRAY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0.GSR.OR_1675  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0.GSR.OR_1676  (
    .I0(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_SFD_ENABLE ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_COUNT_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6.GSR.OR_1677  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG1_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1.GSR.OR_1678  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RX_ER_REG1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1.GSR.OR_1679  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0.GSR.OR_1680  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WAG_READSYNC_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0.GSR.OR_1681  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1.GSR.OR_1682  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2.GSR.OR_1683  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDRGRAY_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2.GSR.OR_1684  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1.GSR.OR_1685  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6.GSR.OR_1686  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_IFG_CNTR_6.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT.GSR.OR_1687  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3.GSR.OR_1688  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1.GSR.OR_1689  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT.GSR.OR_1690  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3.GSR.OR_1691  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1.GSR.OR_1692  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT.GSR.OR_1693  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3.GSR.OR_1694  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1.GSR.OR_1695  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0.GSR.OR_1696  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_RAG_WRITESYNC_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT.GSR.OR_1697  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_RESET_OUT.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3.GSR.OR_1698  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R3.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0.GSR.OR_1699  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_RD_ADDR_0.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2.GSR.OR_1700  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_TX_RESET_I_R2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2.GSR.OR_1701  (
    .I0(\BU2/U0/TRIMAC_INST_INT_TX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_R2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2.GSR.OR_1702  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_RX_RESET_I_R2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1.GSR.OR_1703  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_WR_ADDR_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2.GSR.OR_1704  (
    .I0(\BU2/U0/TRIMAC_INST_INT_RX_RST_ASYNCH ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_R2.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5.GSR.OR_1705  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_TX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_TX_GEN_GMII_TXD_TO_PHY_5.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1.GSR.OR_1706  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_GMII_MII_RX_GEN_RXD_REG4_1.GSR.OR )
  );
  X_OR2 \BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2.GSR.OR_1707  (
    .I0(\BU2/U0/TRIMAC_INST_SYNC_GMII_MII_RX_RESET_I_RESET_OUT ),
    .I1(GSR),
    .O(\BU2/U0/TRIMAC_INST_RXGEN_RX_FIFO_NEXT_WR_ADDR_2.GSR.OR )
  );
  X_ZERO NlwBlock_temac1_GND (
    .O(GND)
  );
  X_ONE NlwBlock_temac1_VCC (
    .O(VCC)
  );
endmodule

