library verilog;
use verilog.vl_types.all;
entity frame_typ is
end frame_typ;
