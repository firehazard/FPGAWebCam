library verilog;
use verilog.vl_types.all;
entity testbench is
    generic(
        dly             : integer := 6000
    );
end testbench;
