library verilog;
use verilog.vl_types.all;
entity sccb_testbench is
end sccb_testbench;
